magic
tech sky130A
magscale 1 2
timestamp 1754964561
<< metal1 >>
rect 7104 27983 7433 27985
rect 6226 27582 6236 27983
rect 7095 27582 7433 27983
rect 21013 2035 21023 2403
rect 21328 2035 21338 2403
<< via1 >>
rect 6236 27582 7095 27983
rect 21023 2035 21328 2403
<< metal2 >>
rect 2046 30457 2446 30467
rect 2046 30047 2446 30057
rect 10489 30171 10889 30362
rect 25088 30171 25439 30181
rect 10489 29859 25088 30171
rect 25088 29849 25439 29859
rect 11068 29793 11226 29803
rect 11068 29294 11226 29599
rect 4796 29136 11226 29294
rect 4796 14947 4954 29136
rect 6236 27983 7095 27993
rect 6236 27572 7095 27582
rect 5273 19462 5373 19472
rect 5373 19410 5977 19462
rect 5273 19375 5373 19385
rect 4796 14875 8161 14947
rect 4796 12094 4954 14875
rect 21526 14480 22053 14481
rect 21513 14474 22053 14480
rect 21513 14471 22054 14474
rect 21513 13979 21526 14471
rect 22053 14464 22054 14471
rect 22053 13979 22054 13980
rect 21526 13970 22054 13979
rect 21526 13969 22053 13970
rect 9591 13059 10125 13069
rect 9591 12815 10125 12927
rect 12349 12101 12894 12111
rect 4796 12022 7759 12094
rect 5273 11125 5373 11135
rect 5373 11053 5749 11125
rect 12349 11092 12894 11926
rect 13324 11262 20778 11398
rect 5273 11043 5373 11053
rect 13324 10349 13473 11262
rect 12919 10295 13473 10349
rect 13324 10293 13473 10295
rect 11366 10242 11466 10252
rect 11466 10172 11840 10226
rect 11366 10162 11466 10172
rect 4365 9919 4498 9929
rect 4498 9818 5684 9919
rect 4365 9808 4498 9818
rect 3925 9768 4058 9778
rect 4058 9668 5676 9768
rect 20642 9686 20778 11262
rect 3925 9658 4058 9668
rect 20487 9550 20778 9686
rect 11237 8566 11709 9222
rect 4528 8529 4703 8539
rect 4703 8129 5360 8529
rect 4528 8119 4703 8129
rect 10766 8094 11709 8566
rect 26466 8168 26867 8178
rect 26466 7607 26867 7617
rect 27234 5535 27414 5545
rect 26879 5380 27234 5535
rect 27234 5370 27414 5380
rect 13750 2396 16043 2406
rect 13750 2171 16043 2181
rect 21023 2403 21328 2413
rect 11778 678 11958 688
rect 18082 678 18134 2106
rect 11768 626 11778 678
rect 11958 626 18134 678
rect 11778 601 11958 611
rect 15642 455 15822 465
rect 18408 455 18460 2115
rect 18704 2087 18794 2097
rect 21023 2025 21328 2035
rect 18704 1908 18794 1988
rect 18704 1836 21155 1908
rect 19506 839 19687 1836
rect 24343 1577 24475 1587
rect 24343 1418 24475 1428
rect 19506 680 19687 690
rect 15822 403 18460 455
rect 15642 385 15822 395
<< via2 >>
rect 2046 30057 2446 30457
rect 25088 29859 25439 30171
rect 11068 29599 11226 29793
rect 6236 27582 7095 27983
rect 5273 19385 5373 19462
rect 21526 14464 22053 14471
rect 21526 13980 22054 14464
rect 21526 13979 22053 13980
rect 9591 12927 10125 13059
rect 12349 11926 12894 12101
rect 5273 11053 5373 11125
rect 11366 10172 11466 10242
rect 4365 9818 4498 9919
rect 3925 9668 4058 9768
rect 4528 8129 4703 8529
rect 26466 7617 26867 8168
rect 27234 5380 27414 5535
rect 13750 2181 16043 2396
rect 11778 611 11958 678
rect 18704 1988 18794 2087
rect 21023 2035 21328 2403
rect 24343 1428 24475 1577
rect 19506 690 19687 839
rect 15642 395 15822 455
<< metal3 >>
rect 2036 30457 2456 30462
rect 2036 30057 2046 30457
rect 2446 30057 2456 30457
rect 2036 30052 2456 30057
rect 25078 30171 25449 30176
rect 2769 13560 2869 29931
rect 25078 29859 25088 30171
rect 25439 29859 25449 30171
rect 25078 29854 25449 29859
rect 11058 29793 11236 29798
rect 11058 29599 11068 29793
rect 11226 29599 11236 29793
rect 11058 29594 11236 29599
rect 6226 27983 7105 27988
rect 6226 27582 6236 27983
rect 7095 27582 7105 27983
rect 6226 27577 7105 27582
rect 5490 24045 5500 24115
rect 5598 24045 5683 24115
rect 5263 19462 5383 19467
rect 5263 19385 5273 19462
rect 5373 19385 5383 19462
rect 5263 19380 5383 19385
rect 21516 14471 22063 14476
rect 21516 13979 21526 14471
rect 22053 14469 22063 14471
rect 22053 14464 22064 14469
rect 22054 13980 22064 14464
rect 22053 13979 22064 13980
rect 21516 13975 22064 13979
rect 21516 13974 22063 13975
rect 2769 13460 11466 13560
rect 9581 13059 10135 13064
rect 9581 12927 9591 13059
rect 10125 12927 10135 13059
rect 9581 12922 10135 12927
rect 5263 11125 5383 11130
rect 5263 11053 5273 11125
rect 5373 11053 5383 11125
rect 5263 11048 5383 11053
rect 11366 10247 11466 13460
rect 12339 12101 12904 12106
rect 12339 11926 12349 12101
rect 12894 11926 12904 12101
rect 12339 11921 12904 11926
rect 11356 10242 11476 10247
rect 11356 10172 11366 10242
rect 11466 10172 11476 10242
rect 11356 10167 11476 10172
rect 4355 9919 4508 9924
rect 4355 9818 4365 9919
rect 4498 9818 4508 9919
rect 4355 9813 4508 9818
rect 3915 9768 4068 9773
rect 3915 9668 3925 9768
rect 4058 9668 4068 9768
rect 3915 9663 4068 9668
rect 4518 8529 4713 8534
rect 2862 8129 2868 8529
rect 3266 8129 4528 8529
rect 4703 8129 4713 8529
rect 4518 8124 4713 8129
rect 5482 2402 5847 2407
rect 2985 2035 2991 2402
rect 3356 2401 5848 2402
rect 3356 2036 5482 2401
rect 5847 2036 5848 2401
rect 3356 2035 5848 2036
rect 5482 2030 5847 2035
rect 12025 1365 12113 9138
rect 13137 8729 13225 9108
rect 13127 8634 13137 8729
rect 13225 8634 13235 8729
rect 26456 8168 26877 8173
rect 26456 7617 26466 8168
rect 26867 7617 26877 8168
rect 26456 7612 26877 7617
rect 27224 5535 27424 5540
rect 27224 5380 27234 5535
rect 27414 5380 27424 5535
rect 27224 5375 27424 5380
rect 20726 3860 21115 4017
rect 13740 2396 16053 2401
rect 13740 2181 13750 2396
rect 16043 2181 16053 2396
rect 13740 2176 16053 2181
rect 18694 2087 18804 2092
rect 18694 1988 18704 2087
rect 18794 1988 18804 2087
rect 18694 1983 18804 1988
rect 7914 1185 12113 1365
rect 7914 785 8094 1185
rect 19496 839 19697 844
rect 7904 620 7914 785
rect 8094 620 8104 785
rect 19496 690 19506 839
rect 19687 690 19697 839
rect 19496 685 19697 690
rect 20726 841 20883 3860
rect 21013 2403 21338 2408
rect 21013 2035 21023 2403
rect 21328 2035 21338 2403
rect 21013 2030 21338 2035
rect 24333 1577 24485 1582
rect 24333 1428 24343 1577
rect 24475 1428 24485 1577
rect 24333 1423 24485 1428
rect 20726 684 23370 841
rect 23550 684 23556 841
rect 11768 678 11968 683
rect 11768 601 11778 678
rect 11958 601 11968 678
rect 15632 455 15832 460
rect 15632 385 15642 455
rect 15822 385 15832 455
<< via3 >>
rect 2046 30057 2446 30457
rect 25088 29859 25439 30171
rect 11068 29599 11226 29793
rect 6236 27582 7095 27983
rect 5500 24045 5598 24115
rect 5273 19385 5373 19462
rect 21526 14464 22053 14471
rect 21526 13980 22054 14464
rect 21526 13979 22053 13980
rect 9591 12927 10125 13059
rect 5273 11053 5373 11125
rect 12349 11926 12894 12101
rect 4365 9818 4498 9919
rect 3925 9668 4058 9768
rect 2868 8129 3266 8529
rect 2991 2035 3356 2402
rect 5482 2036 5847 2401
rect 13137 8634 13225 8729
rect 26466 7617 26867 8168
rect 27234 5380 27414 5535
rect 13750 2181 16043 2396
rect 7914 620 8094 785
rect 19506 690 19687 839
rect 21023 2035 21328 2403
rect 24343 1428 24475 1577
rect 23370 684 23550 841
rect 11778 611 11958 678
rect 11778 601 11958 611
rect 15642 395 15822 455
rect 15642 385 15822 395
<< metal4 >>
rect 200 1000 600 44152
rect 800 43931 1200 44152
rect 3006 43931 3066 45152
rect 3558 43931 3618 45152
rect 4110 43931 4170 45152
rect 4662 43931 4722 45152
rect 5214 43931 5274 45152
rect 5766 43931 5826 45152
rect 6318 43931 6378 45152
rect 6870 43931 6930 45152
rect 7422 43931 7482 45152
rect 7974 43931 8034 45152
rect 8526 43931 8586 45152
rect 9078 43931 9138 45152
rect 9630 43931 9690 45152
rect 10182 43931 10242 45152
rect 10734 43931 10794 45152
rect 11286 43931 11346 45152
rect 11838 43931 11898 45152
rect 12390 43931 12450 45152
rect 12942 43931 13002 45152
rect 13494 43931 13554 45152
rect 14046 43931 14106 45152
rect 14598 43931 14658 45152
rect 15150 43931 15210 45152
rect 15702 45058 15762 45152
rect 15702 43931 15763 45058
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 800 43741 15765 43931
rect 800 30457 1200 43741
rect 15702 43740 15763 43741
rect 2045 30457 2447 30458
rect 800 30057 2046 30457
rect 2446 30057 2447 30457
rect 800 27982 1200 30057
rect 2045 30056 2447 30057
rect 11068 29794 11226 30524
rect 25087 30171 25440 30172
rect 28400 30171 28800 44152
rect 25087 29859 25088 30171
rect 25439 29859 28800 30171
rect 25087 29858 25440 29859
rect 11067 29793 11227 29794
rect 11067 29599 11068 29793
rect 11226 29599 11227 29793
rect 11067 29598 11227 29599
rect 6235 27983 7096 27984
rect 6235 27982 6236 27983
rect 800 27582 6236 27982
rect 7095 27582 7096 27983
rect 800 8529 1200 27582
rect 6235 27581 7096 27582
rect 5499 24115 5599 24116
rect 4365 24045 5500 24115
rect 5598 24045 5642 24115
rect 4365 9920 4498 24045
rect 5499 24044 5599 24045
rect 5272 19462 5374 19463
rect 5272 19385 5273 19462
rect 5373 19385 5374 19462
rect 5272 19384 5374 19385
rect 5273 11126 5373 19384
rect 9591 14471 22127 14474
rect 9591 13981 21526 14471
rect 22053 14464 22127 14471
rect 28400 14464 28800 29859
rect 9591 13060 10125 13981
rect 12077 13974 12894 13981
rect 21525 13979 21526 13981
rect 22054 13981 28800 14464
rect 22054 13980 22055 13981
rect 22053 13979 22055 13980
rect 21525 13978 22054 13979
rect 9590 13059 10126 13060
rect 9590 12927 9591 13059
rect 10125 12927 10126 13059
rect 9590 12926 10126 12927
rect 12349 12102 12894 13974
rect 12348 12101 12895 12102
rect 12348 11926 12349 12101
rect 12894 11926 12895 12101
rect 12348 11925 12895 11926
rect 5272 11125 5374 11126
rect 5272 11053 5273 11125
rect 5373 11053 5374 11125
rect 5272 11052 5374 11053
rect 4364 9919 4499 9920
rect 4364 9818 4365 9919
rect 4498 9818 4499 9919
rect 4364 9817 4499 9818
rect 3924 9768 4059 9769
rect 3924 9668 3925 9768
rect 4058 9668 4059 9768
rect 3924 9667 4059 9668
rect 2867 8529 3267 8530
rect 800 8129 2868 8529
rect 3266 8129 3267 8529
rect 800 2402 1200 8129
rect 2867 8128 3267 8129
rect 2990 2402 3357 2403
rect 800 2035 2991 2402
rect 3356 2035 3357 2402
rect 800 1000 1200 2035
rect 2990 2034 3357 2035
rect 3925 1561 4058 9667
rect 13136 8729 13226 8730
rect 10886 8634 13137 8729
rect 13225 8634 13226 8729
rect 13136 8633 13226 8634
rect 26465 8168 26868 8169
rect 28400 8168 28800 13981
rect 26465 7617 26466 8168
rect 26867 7617 28800 8168
rect 26465 7616 26868 7617
rect 27233 5535 27415 5536
rect 27233 5380 27234 5535
rect 27414 5380 27415 5535
rect 27233 5379 27415 5380
rect 21022 2403 21329 2404
rect 21022 2402 21023 2403
rect 5481 2401 21023 2402
rect 5481 2036 5482 2401
rect 5847 2396 21023 2401
rect 5847 2181 13750 2396
rect 16043 2181 21023 2396
rect 5847 2036 21023 2181
rect 5481 2035 21023 2036
rect 21328 2402 21329 2403
rect 21328 2035 21335 2402
rect 21022 2034 21329 2035
rect 24342 1577 24476 1578
rect 24342 1561 24343 1577
rect 3925 1428 24343 1561
rect 24475 1428 24476 1577
rect 24342 1427 24476 1428
rect 24343 1418 24476 1427
rect 19506 840 19687 903
rect 23369 841 23551 842
rect 19505 839 19688 840
rect 7913 785 8095 786
rect 7913 620 7914 785
rect 8094 620 8095 785
rect 19505 690 19506 839
rect 19687 690 19688 839
rect 19505 689 19688 690
rect 7913 619 8095 620
rect 11777 678 11959 679
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 619
rect 11777 601 11778 678
rect 11958 601 11959 678
rect 11777 600 11959 601
rect 11778 0 11958 600
rect 15641 455 15823 456
rect 15641 385 15642 455
rect 15822 385 15823 455
rect 15641 384 15823 385
rect 15642 0 15822 384
rect 19506 188 19687 689
rect 23369 684 23370 841
rect 23550 684 23551 841
rect 23369 683 23551 684
rect 19506 0 19686 188
rect 23370 0 23550 683
rect 27234 0 27414 5379
rect 28400 1000 28800 7617
use BIAS_1  BIAS_1_0 ~/Dalin/X51/magic/bias
timestamp 1754956152
transform -1 0 61672 0 -1 37488
box 33736 9131 56010 23507
use COMP_2  COMP_2_0 ~/Dalin/X51/magic/COMP
timestamp 1754963760
transform 1 0 -5506 0 1 12999
box 10603 -7294 16407 -165
use delay_1  delay_1_0 ~/Dalin/X51/magic/slowsw
timestamp 1754019877
transform 1 0 -33625 0 1 30371
box 35948 -1101 58337 12413
use latch_sch  latch_sch_0 ~/Dalin/X51/magic/latch
timestamp 1754960833
transform 1 0 9856 0 1 10939
box 1372 -1870 3610 189
use Timming  Timming_0 ~/Dalin/X51/magic/timming_magic
timestamp 1751928886
transform 1 0 7900 0 1 5005
box 5707 -2926 12653 6071
use VCR  VCR_0 ~/Dalin/X51/magic/VCR
timestamp 1752032521
transform 1 0 20794 0 1 4246
box 309 -2692 6139 3934
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 28400 1000 28800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
