VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_asic
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_asic ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.860000 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 180.000000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 50.000000 ;
    ANTENNADIFFAREA 0.290000 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 30.000000 ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 30.000000 ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.000000 ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.560089 ;
    ANTENNADIFFAREA 781.075195 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 142.000 5.000 144.000 220.760 ;
    END
  END VAPWR
  OBS
      LAYER pwell ;
        RECT 13.100 150.910 28.430 212.020 ;
      LAYER nwell ;
        RECT 30.105 152.105 54.315 156.075 ;
      LAYER pwell ;
        RECT 37.100 135.470 67.210 141.395 ;
        RECT 36.850 134.915 67.210 135.470 ;
        RECT 37.100 123.105 67.210 134.915 ;
        RECT 68.105 140.675 88.245 141.440 ;
        RECT 68.105 135.505 68.870 140.675 ;
        RECT 74.040 135.505 75.590 140.675 ;
        RECT 80.760 135.505 82.310 140.675 ;
        RECT 87.480 135.505 88.245 140.675 ;
        RECT 68.105 133.955 88.245 135.505 ;
        RECT 68.105 128.785 68.870 133.955 ;
        RECT 74.040 128.785 75.590 133.955 ;
        RECT 80.760 128.785 82.310 133.955 ;
        RECT 87.480 128.785 88.245 133.955 ;
        RECT 68.105 127.235 88.245 128.785 ;
        RECT 68.105 122.065 68.870 127.235 ;
        RECT 74.040 122.065 75.590 127.235 ;
        RECT 80.760 122.065 82.310 127.235 ;
        RECT 87.480 122.065 88.245 127.235 ;
        RECT 54.065 121.420 54.535 121.735 ;
        RECT 29.470 99.140 54.535 121.420 ;
        RECT 68.105 121.300 88.245 122.065 ;
        RECT 78.075 117.385 100.355 119.385 ;
        RECT 55.795 111.805 100.355 117.385 ;
        RECT 55.830 105.445 100.355 111.025 ;
        RECT 55.830 103.445 78.110 105.445 ;
        RECT 54.065 98.595 54.535 99.140 ;
      LAYER nwell ;
        RECT 30.730 83.770 53.310 96.740 ;
        RECT 40.780 71.750 53.310 75.720 ;
        RECT 56.170 71.750 100.380 96.740 ;
        RECT 103.010 72.320 109.000 94.900 ;
        RECT 39.305 59.285 51.935 63.100 ;
        RECT 29.305 59.130 51.935 59.285 ;
        RECT 29.305 54.445 51.885 59.130 ;
        RECT 59.235 55.425 64.415 55.575 ;
        RECT 29.305 54.315 53.835 54.445 ;
        RECT 29.865 43.675 39.525 54.315 ;
        RECT 44.195 43.550 53.835 54.315 ;
        RECT 59.180 52.110 64.575 55.425 ;
        RECT 59.235 52.035 64.415 52.110 ;
      LAYER pwell ;
        RECT 56.175 45.960 67.295 49.540 ;
        RECT 26.415 28.965 42.975 43.285 ;
        RECT 44.345 39.705 48.825 43.285 ;
        RECT 49.205 39.710 53.685 43.290 ;
        RECT 69.655 12.205 82.025 54.315 ;
        RECT 82.135 37.150 101.505 49.730 ;
        RECT 82.115 24.515 91.555 36.795 ;
        RECT 82.115 12.205 91.555 24.485 ;
        RECT 92.740 12.205 99.190 32.025 ;
        RECT 107.395 18.105 119.975 40.635 ;
      LAYER nwell ;
        RECT 122.670 37.255 129.640 40.785 ;
        RECT 122.670 24.645 134.140 37.255 ;
      LAYER pwell ;
        RECT 106.320 8.345 121.210 15.925 ;
        RECT 122.040 8.815 134.620 20.095 ;
      LAYER li1 ;
        RECT 12.025 213.100 28.970 213.110 ;
        RECT 12.025 211.555 29.205 213.100 ;
        RECT 12.025 181.550 13.580 211.555 ;
        RECT 13.930 209.030 14.280 211.190 ;
        RECT 13.930 182.030 14.280 184.190 ;
        RECT 14.760 181.550 14.930 211.555 ;
        RECT 15.410 209.030 15.760 211.190 ;
        RECT 15.410 182.030 15.760 184.190 ;
        RECT 16.240 181.550 16.410 211.555 ;
        RECT 16.890 209.030 17.240 211.190 ;
        RECT 16.890 182.030 17.240 184.190 ;
        RECT 17.720 181.550 17.890 211.555 ;
        RECT 18.370 209.030 18.720 211.190 ;
        RECT 18.370 182.030 18.720 184.190 ;
        RECT 19.200 181.550 19.370 211.555 ;
        RECT 19.850 209.030 20.200 211.190 ;
        RECT 19.850 182.030 20.200 184.190 ;
        RECT 20.680 181.550 20.850 211.555 ;
        RECT 21.330 209.030 21.680 211.190 ;
        RECT 21.330 182.030 21.680 184.190 ;
        RECT 22.160 181.550 22.330 211.555 ;
        RECT 22.810 209.030 23.160 211.190 ;
        RECT 22.810 182.030 23.160 184.190 ;
        RECT 23.640 181.550 23.810 211.555 ;
        RECT 24.290 209.030 24.640 211.190 ;
        RECT 24.290 182.030 24.640 184.190 ;
        RECT 25.120 181.550 25.290 211.555 ;
        RECT 25.770 209.030 26.120 211.190 ;
        RECT 25.770 182.030 26.120 184.190 ;
        RECT 26.600 181.550 26.770 211.555 ;
        RECT 27.250 209.030 27.600 211.190 ;
        RECT 27.250 182.030 27.600 184.190 ;
        RECT 27.950 181.550 29.205 211.555 ;
        RECT 12.025 181.380 29.205 181.550 ;
        RECT 12.025 151.470 13.580 181.380 ;
        RECT 13.930 178.740 14.280 180.900 ;
        RECT 13.930 151.740 14.280 153.900 ;
        RECT 14.760 151.470 14.930 181.380 ;
        RECT 15.410 178.740 15.760 180.900 ;
        RECT 15.410 151.740 15.760 153.900 ;
        RECT 16.240 151.470 16.410 181.380 ;
        RECT 16.890 178.740 17.240 180.900 ;
        RECT 16.890 151.740 17.240 153.900 ;
        RECT 17.720 151.470 17.890 181.380 ;
        RECT 18.370 178.740 18.720 180.900 ;
        RECT 18.370 151.740 18.720 153.900 ;
        RECT 19.200 151.470 19.370 181.380 ;
        RECT 19.850 178.740 20.200 180.900 ;
        RECT 19.850 151.740 20.200 153.900 ;
        RECT 20.680 151.470 20.850 181.380 ;
        RECT 21.330 178.740 21.680 180.900 ;
        RECT 21.330 151.740 21.680 153.900 ;
        RECT 22.160 151.470 22.330 181.380 ;
        RECT 22.810 178.740 23.160 180.900 ;
        RECT 22.810 151.740 23.160 153.900 ;
        RECT 23.640 151.470 23.810 181.380 ;
        RECT 24.290 178.740 24.640 180.900 ;
        RECT 24.290 151.740 24.640 153.900 ;
        RECT 25.120 151.470 25.290 181.380 ;
        RECT 25.770 178.740 26.120 180.900 ;
        RECT 25.770 151.740 26.120 153.900 ;
        RECT 26.600 151.470 26.770 181.380 ;
        RECT 27.250 178.740 27.600 180.900 ;
        RECT 27.250 151.740 27.600 153.900 ;
        RECT 27.950 151.470 29.205 181.380 ;
        RECT 30.160 156.420 54.415 156.515 ;
        RECT 30.110 155.490 54.520 156.420 ;
        RECT 30.110 152.735 30.800 155.490 ;
        RECT 31.395 154.825 41.395 154.995 ;
        RECT 31.165 153.570 31.335 154.610 ;
        RECT 41.455 153.570 41.625 154.610 ;
        RECT 31.395 153.185 41.395 153.355 ;
        RECT 42.125 152.735 42.295 155.490 ;
        RECT 43.025 154.825 53.025 154.995 ;
        RECT 42.795 153.570 42.965 154.610 ;
        RECT 53.085 153.570 53.255 154.610 ;
        RECT 43.025 153.185 53.025 153.355 ;
        RECT 53.740 152.735 54.520 155.490 ;
        RECT 30.110 151.675 54.520 152.735 ;
        RECT 12.025 150.140 29.205 151.470 ;
        RECT 36.675 140.915 88.165 141.785 ;
        RECT 36.675 139.870 37.475 140.915 ;
        RECT 37.930 140.215 40.090 140.565 ;
        RECT 49.430 140.215 51.590 140.565 ;
        RECT 51.885 139.870 52.375 140.915 ;
        RECT 52.720 140.215 54.880 140.565 ;
        RECT 64.220 140.215 66.380 140.565 ;
        RECT 66.850 140.135 88.165 140.915 ;
        RECT 66.850 139.870 69.410 140.135 ;
        RECT 36.675 139.315 69.410 139.870 ;
        RECT 36.675 138.405 37.475 139.315 ;
        RECT 37.930 138.735 40.090 139.085 ;
        RECT 49.430 138.735 51.590 139.085 ;
        RECT 51.885 138.405 52.375 139.315 ;
        RECT 52.720 138.735 54.880 139.085 ;
        RECT 64.220 138.735 66.380 139.085 ;
        RECT 66.850 138.405 69.410 139.315 ;
        RECT 36.675 137.850 69.410 138.405 ;
        RECT 36.675 136.935 37.475 137.850 ;
        RECT 37.930 137.255 40.090 137.605 ;
        RECT 49.430 137.255 51.590 137.605 ;
        RECT 51.885 136.935 52.375 137.850 ;
        RECT 52.720 137.255 54.880 137.605 ;
        RECT 64.220 137.255 66.380 137.605 ;
        RECT 66.850 136.935 69.410 137.850 ;
        RECT 36.675 136.380 69.410 136.935 ;
        RECT 36.675 135.470 37.475 136.380 ;
        RECT 37.930 135.775 40.090 136.125 ;
        RECT 49.430 135.775 51.590 136.125 ;
        RECT 51.885 135.470 52.375 136.380 ;
        RECT 52.720 135.775 54.880 136.125 ;
        RECT 64.220 135.775 66.380 136.125 ;
        RECT 66.850 136.045 69.410 136.380 ;
        RECT 69.720 136.355 73.190 139.825 ;
        RECT 73.500 136.045 76.130 140.135 ;
        RECT 76.440 136.355 79.910 139.825 ;
        RECT 80.220 136.045 82.850 140.135 ;
        RECT 83.160 136.355 86.630 139.825 ;
        RECT 86.940 136.045 88.165 140.135 ;
        RECT 66.850 135.470 88.165 136.045 ;
        RECT 36.675 134.915 88.165 135.470 ;
        RECT 36.675 134.005 37.475 134.915 ;
        RECT 37.930 134.295 40.090 134.645 ;
        RECT 49.430 134.295 51.590 134.645 ;
        RECT 51.885 134.005 52.375 134.915 ;
        RECT 52.720 134.295 54.880 134.645 ;
        RECT 64.220 134.295 66.380 134.645 ;
        RECT 66.850 134.095 88.165 134.915 ;
        RECT 66.850 134.005 69.270 134.095 ;
        RECT 36.675 133.775 69.270 134.005 ;
        RECT 73.585 133.775 76.000 134.095 ;
        RECT 80.365 133.775 82.665 134.095 ;
        RECT 87.080 133.775 88.165 134.095 ;
        RECT 36.675 133.450 88.165 133.775 ;
        RECT 36.675 132.540 37.475 133.450 ;
        RECT 37.930 132.815 40.090 133.165 ;
        RECT 49.430 132.815 51.590 133.165 ;
        RECT 51.885 132.540 52.375 133.450 ;
        RECT 66.850 133.415 88.165 133.450 ;
        RECT 52.720 132.815 54.880 133.165 ;
        RECT 64.220 132.815 66.380 133.165 ;
        RECT 66.850 132.540 69.410 133.415 ;
        RECT 36.675 131.985 69.410 132.540 ;
        RECT 36.675 131.040 37.475 131.985 ;
        RECT 37.930 131.335 40.090 131.685 ;
        RECT 49.430 131.335 51.590 131.685 ;
        RECT 51.885 131.040 52.375 131.985 ;
        RECT 52.720 131.335 54.880 131.685 ;
        RECT 64.220 131.335 66.380 131.685 ;
        RECT 66.850 131.040 69.410 131.985 ;
        RECT 36.675 130.485 69.410 131.040 ;
        RECT 36.675 129.505 37.475 130.485 ;
        RECT 37.930 129.855 40.090 130.205 ;
        RECT 49.430 129.855 51.590 130.205 ;
        RECT 51.885 129.505 52.375 130.485 ;
        RECT 52.720 129.855 54.880 130.205 ;
        RECT 64.220 129.855 66.380 130.205 ;
        RECT 66.850 129.505 69.410 130.485 ;
        RECT 69.720 129.635 73.190 133.105 ;
        RECT 36.675 129.325 69.410 129.505 ;
        RECT 73.500 129.325 76.130 133.415 ;
        RECT 76.440 129.635 79.910 133.105 ;
        RECT 80.220 129.325 82.850 133.415 ;
        RECT 83.160 129.635 86.630 133.105 ;
        RECT 86.940 129.325 88.165 133.415 ;
        RECT 36.675 128.950 88.165 129.325 ;
        RECT 36.675 128.075 37.475 128.950 ;
        RECT 37.930 128.375 40.090 128.725 ;
        RECT 49.430 128.375 51.590 128.725 ;
        RECT 51.885 128.075 52.375 128.950 ;
        RECT 52.720 128.375 54.880 128.725 ;
        RECT 64.220 128.375 66.380 128.725 ;
        RECT 66.850 128.075 88.165 128.950 ;
        RECT 36.675 127.520 88.165 128.075 ;
        RECT 36.675 126.610 37.475 127.520 ;
        RECT 37.930 126.895 40.090 127.245 ;
        RECT 49.430 126.895 51.590 127.245 ;
        RECT 51.885 126.610 52.375 127.520 ;
        RECT 52.720 126.895 54.880 127.245 ;
        RECT 64.220 126.895 66.380 127.245 ;
        RECT 66.850 126.695 88.165 127.520 ;
        RECT 66.850 126.610 69.410 126.695 ;
        RECT 36.675 126.055 69.410 126.610 ;
        RECT 36.675 125.075 37.475 126.055 ;
        RECT 37.930 125.415 40.090 125.765 ;
        RECT 49.430 125.415 51.590 125.765 ;
        RECT 51.885 125.075 52.375 126.055 ;
        RECT 52.720 125.415 54.880 125.765 ;
        RECT 64.220 125.415 66.380 125.765 ;
        RECT 66.850 125.075 69.410 126.055 ;
        RECT 36.675 124.520 69.410 125.075 ;
        RECT 36.675 123.505 37.475 124.520 ;
        RECT 37.930 123.935 40.090 124.285 ;
        RECT 49.430 123.935 51.590 124.285 ;
        RECT 51.885 123.505 52.375 124.520 ;
        RECT 52.720 123.935 54.880 124.285 ;
        RECT 64.220 123.935 66.380 124.285 ;
        RECT 66.850 123.505 69.410 124.520 ;
        RECT 36.675 123.450 69.410 123.505 ;
        RECT 28.710 122.605 69.410 123.450 ;
        RECT 69.720 122.915 73.190 126.385 ;
        RECT 73.500 122.605 76.130 126.695 ;
        RECT 76.440 122.915 79.910 126.385 ;
        RECT 80.220 122.605 82.850 126.695 ;
        RECT 83.160 122.915 86.630 126.385 ;
        RECT 86.940 122.605 88.165 126.695 ;
        RECT 28.710 120.840 88.165 122.605 ;
        RECT 28.710 99.770 29.905 120.840 ;
        RECT 30.740 120.340 31.280 120.510 ;
        RECT 30.400 100.280 30.570 120.280 ;
        RECT 31.450 100.280 31.620 120.280 ;
        RECT 30.740 100.050 31.280 100.220 ;
        RECT 32.140 99.770 32.310 120.840 ;
        RECT 33.170 120.340 33.710 120.510 ;
        RECT 32.830 100.280 33.000 120.280 ;
        RECT 33.880 100.280 34.050 120.280 ;
        RECT 33.170 100.050 33.710 100.220 ;
        RECT 34.570 99.770 34.740 120.840 ;
        RECT 35.600 120.340 36.140 120.510 ;
        RECT 35.260 100.280 35.430 120.280 ;
        RECT 36.310 100.280 36.480 120.280 ;
        RECT 35.600 100.050 36.140 100.220 ;
        RECT 37.000 99.770 37.170 120.840 ;
        RECT 38.030 120.340 38.570 120.510 ;
        RECT 37.690 100.280 37.860 120.280 ;
        RECT 38.740 100.280 38.910 120.280 ;
        RECT 38.030 100.050 38.570 100.220 ;
        RECT 39.430 99.770 39.600 120.840 ;
        RECT 40.460 120.340 41.000 120.510 ;
        RECT 40.120 100.280 40.290 120.280 ;
        RECT 41.170 100.280 41.340 120.280 ;
        RECT 40.460 100.050 41.000 100.220 ;
        RECT 41.860 99.770 42.030 120.840 ;
        RECT 42.890 120.340 43.430 120.510 ;
        RECT 42.550 100.280 42.720 120.280 ;
        RECT 43.600 100.280 43.770 120.280 ;
        RECT 42.890 100.050 43.430 100.220 ;
        RECT 44.290 99.770 44.460 120.840 ;
        RECT 45.320 120.340 45.860 120.510 ;
        RECT 44.980 100.280 45.150 120.280 ;
        RECT 46.030 100.280 46.200 120.280 ;
        RECT 45.320 100.050 45.860 100.220 ;
        RECT 46.720 99.770 46.890 120.840 ;
        RECT 47.750 120.340 48.290 120.510 ;
        RECT 47.410 100.280 47.580 120.280 ;
        RECT 48.460 100.280 48.630 120.280 ;
        RECT 47.750 100.050 48.290 100.220 ;
        RECT 49.150 99.770 49.320 120.840 ;
        RECT 50.180 120.340 50.720 120.510 ;
        RECT 49.840 100.280 50.010 120.280 ;
        RECT 50.890 100.280 51.060 120.280 ;
        RECT 50.180 100.050 50.720 100.220 ;
        RECT 51.580 99.770 51.750 120.840 ;
        RECT 52.610 120.340 53.150 120.510 ;
        RECT 53.815 120.340 88.165 120.840 ;
        RECT 52.270 100.280 52.440 120.280 ;
        RECT 53.320 100.280 53.490 120.280 ;
        RECT 53.815 118.880 100.775 120.340 ;
        RECT 53.815 116.820 78.580 118.880 ;
        RECT 79.215 118.285 99.215 118.455 ;
        RECT 53.815 112.285 56.260 116.820 ;
        RECT 56.935 116.285 76.935 116.455 ;
        RECT 56.705 113.075 56.875 116.115 ;
        RECT 76.995 113.075 77.165 116.115 ;
        RECT 56.935 112.735 76.935 112.905 ;
        RECT 77.630 112.285 78.580 116.820 ;
        RECT 78.985 113.075 79.155 118.115 ;
        RECT 99.275 113.075 99.445 118.115 ;
        RECT 79.215 112.735 99.215 112.905 ;
        RECT 99.825 112.285 100.775 118.880 ;
        RECT 53.815 110.480 100.775 112.285 ;
        RECT 53.815 103.920 56.305 110.480 ;
        RECT 56.970 109.925 76.970 110.095 ;
        RECT 56.740 104.715 56.910 109.755 ;
        RECT 77.030 104.715 77.200 109.755 ;
        RECT 77.565 105.945 78.550 110.480 ;
        RECT 79.215 109.925 99.215 110.095 ;
        RECT 78.985 106.715 79.155 109.755 ;
        RECT 99.275 106.715 99.445 109.755 ;
        RECT 79.215 106.375 99.215 106.545 ;
        RECT 99.825 105.945 100.775 110.480 ;
        RECT 77.565 105.405 100.775 105.945 ;
        RECT 56.970 104.375 76.970 104.545 ;
        RECT 53.815 103.915 56.315 103.920 ;
        RECT 77.660 103.915 78.000 105.405 ;
        RECT 53.815 103.480 78.015 103.915 ;
        RECT 52.610 100.050 53.150 100.220 ;
        RECT 53.815 99.770 54.470 103.480 ;
        RECT 28.710 98.655 54.470 99.770 ;
        RECT 56.070 96.830 100.540 96.835 ;
        RECT 30.680 95.980 100.540 96.830 ;
        RECT 30.680 95.955 56.820 95.980 ;
        RECT 30.680 90.205 31.345 95.955 ;
        RECT 32.020 95.490 52.020 95.660 ;
        RECT 31.790 93.735 31.960 95.275 ;
        RECT 52.080 93.735 52.250 95.275 ;
        RECT 32.020 93.350 52.020 93.520 ;
        RECT 32.020 92.810 52.020 92.980 ;
        RECT 31.790 91.055 31.960 92.595 ;
        RECT 52.080 91.055 52.250 92.595 ;
        RECT 32.020 90.670 52.020 90.840 ;
        RECT 52.585 90.205 56.820 95.955 ;
        RECT 57.460 95.490 77.460 95.660 ;
        RECT 30.680 89.020 56.820 90.205 ;
        RECT 30.680 84.435 31.345 89.020 ;
        RECT 32.020 88.490 52.020 88.660 ;
        RECT 31.790 85.235 31.960 88.275 ;
        RECT 52.080 85.235 52.250 88.275 ;
        RECT 32.020 84.850 52.020 85.020 ;
        RECT 30.680 84.400 42.745 84.435 ;
        RECT 30.680 84.395 51.935 84.400 ;
        RECT 52.585 84.395 56.820 89.020 ;
        RECT 57.230 85.235 57.400 95.275 ;
        RECT 77.520 85.235 77.690 95.275 ;
        RECT 57.460 84.850 77.460 85.020 ;
        RECT 30.680 84.330 56.820 84.395 ;
        RECT 78.190 84.330 78.360 95.980 ;
        RECT 79.090 95.490 99.090 95.660 ;
        RECT 78.860 85.235 79.030 95.275 ;
        RECT 99.150 85.235 99.320 95.275 ;
        RECT 99.760 94.960 100.510 95.980 ;
        RECT 99.760 94.240 109.155 94.960 ;
        RECT 79.090 84.850 99.090 85.020 ;
        RECT 99.760 84.330 103.685 94.240 ;
        RECT 104.475 93.670 105.015 93.840 ;
        RECT 30.680 84.160 103.685 84.330 ;
        RECT 30.680 83.705 56.820 84.160 ;
        RECT 30.765 83.685 56.820 83.705 ;
        RECT 40.280 75.110 56.820 83.685 ;
        RECT 57.460 83.470 77.460 83.640 ;
        RECT 40.255 75.040 56.820 75.110 ;
        RECT 40.255 72.410 41.345 75.040 ;
        RECT 42.070 74.470 52.020 74.640 ;
        RECT 41.840 73.215 42.010 74.255 ;
        RECT 52.080 73.215 52.250 74.255 ;
        RECT 42.070 72.830 52.020 73.000 ;
        RECT 52.685 72.410 56.820 75.040 ;
        RECT 57.230 73.215 57.400 83.255 ;
        RECT 77.520 73.215 77.690 83.255 ;
        RECT 57.460 72.830 77.460 73.000 ;
        RECT 78.190 72.410 78.360 84.160 ;
        RECT 79.090 83.470 99.090 83.640 ;
        RECT 78.860 73.215 79.030 83.255 ;
        RECT 99.150 73.215 99.320 83.255 ;
        RECT 79.090 72.830 99.090 73.000 ;
        RECT 99.760 72.925 103.685 84.160 ;
        RECT 104.090 73.610 104.260 93.610 ;
        RECT 105.230 73.610 105.400 93.610 ;
        RECT 104.475 73.380 105.015 73.550 ;
        RECT 105.920 72.925 106.090 94.240 ;
        RECT 106.995 93.670 107.535 93.840 ;
        RECT 106.610 73.610 106.780 93.610 ;
        RECT 107.750 73.610 107.920 93.610 ;
        RECT 106.995 73.380 107.535 73.550 ;
        RECT 108.330 72.925 109.155 94.240 ;
        RECT 99.755 72.410 109.155 72.925 ;
        RECT 40.255 70.705 109.155 72.410 ;
        RECT 40.280 70.005 109.155 70.705 ;
        RECT 39.000 64.085 53.890 64.120 ;
        RECT 39.000 64.045 53.955 64.085 ;
        RECT 38.935 62.510 53.955 64.045 ;
        RECT 38.935 59.925 40.130 62.510 ;
        RECT 40.595 61.850 50.645 62.020 ;
        RECT 40.365 60.595 40.535 61.635 ;
        RECT 50.705 60.595 50.875 61.635 ;
        RECT 40.595 60.210 50.645 60.380 ;
        RECT 51.255 59.925 53.955 62.510 ;
        RECT 29.120 58.615 53.955 59.925 ;
        RECT 29.120 55.020 29.980 58.615 ;
        RECT 30.595 58.035 50.595 58.205 ;
        RECT 30.365 55.780 30.535 57.820 ;
        RECT 50.655 55.780 50.825 57.820 ;
        RECT 30.595 55.395 50.595 55.565 ;
        RECT 51.255 55.020 53.955 58.615 ;
        RECT 29.120 53.785 53.955 55.020 ;
        RECT 29.120 49.445 30.545 53.785 ;
        RECT 31.155 53.105 33.555 53.275 ;
        RECT 30.925 50.350 31.095 52.890 ;
        RECT 33.615 50.350 33.785 52.890 ;
        RECT 31.155 49.965 33.555 50.135 ;
        RECT 34.215 49.445 35.225 53.785 ;
        RECT 35.835 53.105 38.235 53.275 ;
        RECT 35.605 50.350 35.775 52.890 ;
        RECT 38.295 50.350 38.465 52.890 ;
        RECT 35.835 49.965 38.235 50.135 ;
        RECT 38.820 49.680 44.890 53.785 ;
        RECT 45.485 53.195 47.885 53.365 ;
        RECT 45.255 50.440 45.425 52.980 ;
        RECT 47.945 50.440 48.115 52.980 ;
        RECT 45.485 50.055 47.885 50.225 ;
        RECT 48.605 49.680 49.525 53.785 ;
        RECT 50.145 53.195 52.545 53.365 ;
        RECT 49.915 50.440 50.085 52.980 ;
        RECT 52.605 50.440 52.775 52.980 ;
        RECT 50.145 50.055 52.545 50.225 ;
        RECT 53.165 49.680 53.955 53.785 ;
        RECT 59.195 54.955 64.590 55.640 ;
        RECT 59.195 52.555 59.970 54.955 ;
        RECT 60.395 54.560 60.895 54.730 ;
        RECT 61.185 54.560 61.685 54.730 ;
        RECT 61.975 54.560 62.475 54.730 ;
        RECT 62.765 54.560 63.265 54.730 ;
        RECT 60.165 53.305 60.335 54.345 ;
        RECT 60.955 53.305 61.125 54.345 ;
        RECT 61.745 53.305 61.915 54.345 ;
        RECT 62.535 53.305 62.705 54.345 ;
        RECT 63.325 53.305 63.495 54.345 ;
        RECT 60.395 52.920 60.895 53.090 ;
        RECT 61.185 52.920 61.685 53.090 ;
        RECT 61.975 52.920 62.475 53.090 ;
        RECT 62.765 52.920 63.265 53.090 ;
        RECT 63.815 52.555 64.590 54.955 ;
        RECT 68.455 53.945 102.225 55.380 ;
        RECT 59.180 51.760 64.590 52.555 ;
        RECT 38.820 49.445 53.955 49.680 ;
        RECT 29.120 49.275 53.955 49.445 ;
        RECT 29.120 48.755 30.545 49.275 ;
        RECT 34.215 48.755 35.225 49.275 ;
        RECT 38.820 48.755 53.955 49.275 ;
        RECT 29.120 48.585 53.955 48.755 ;
        RECT 29.120 44.420 30.545 48.585 ;
        RECT 31.155 47.895 33.555 48.065 ;
        RECT 30.925 45.140 31.095 47.680 ;
        RECT 33.615 45.140 33.785 47.680 ;
        RECT 31.155 44.755 33.555 44.925 ;
        RECT 34.215 44.420 35.225 48.585 ;
        RECT 38.820 48.420 53.955 48.585 ;
        RECT 35.835 47.895 38.235 48.065 ;
        RECT 35.605 45.140 35.775 47.680 ;
        RECT 38.295 45.140 38.465 47.680 ;
        RECT 35.835 44.755 38.235 44.925 ;
        RECT 38.820 44.420 44.890 48.420 ;
        RECT 45.485 47.770 47.885 47.940 ;
        RECT 45.255 45.015 45.425 47.555 ;
        RECT 47.945 45.015 48.115 47.555 ;
        RECT 45.485 44.630 47.885 44.800 ;
        RECT 29.120 44.385 45.075 44.420 ;
        RECT 48.605 44.385 49.525 48.420 ;
        RECT 50.145 47.770 52.545 47.940 ;
        RECT 49.915 45.015 50.085 47.555 ;
        RECT 52.605 45.015 52.775 47.555 ;
        RECT 50.145 44.630 52.545 44.800 ;
        RECT 53.165 44.385 53.955 48.420 ;
        RECT 56.140 49.130 67.330 49.575 ;
        RECT 56.140 46.505 56.645 49.130 ;
        RECT 57.315 48.440 57.815 48.610 ;
        RECT 57.085 47.230 57.255 48.270 ;
        RECT 57.875 47.230 58.045 48.270 ;
        RECT 57.315 46.890 57.815 47.060 ;
        RECT 58.545 46.505 59.365 49.130 ;
        RECT 60.095 48.440 60.595 48.610 ;
        RECT 59.865 47.230 60.035 48.270 ;
        RECT 60.655 47.230 60.825 48.270 ;
        RECT 60.095 46.890 60.595 47.060 ;
        RECT 61.325 46.505 62.145 49.130 ;
        RECT 62.875 48.440 63.375 48.610 ;
        RECT 62.645 47.230 62.815 48.270 ;
        RECT 63.435 47.230 63.605 48.270 ;
        RECT 62.875 46.890 63.375 47.060 ;
        RECT 64.100 46.505 64.925 49.130 ;
        RECT 65.655 48.440 66.155 48.610 ;
        RECT 65.425 47.230 65.595 48.270 ;
        RECT 66.215 47.230 66.385 48.270 ;
        RECT 65.655 46.890 66.155 47.060 ;
        RECT 66.875 46.505 67.330 49.130 ;
        RECT 56.140 45.705 67.330 46.505 ;
        RECT 29.120 43.745 53.955 44.385 ;
        RECT 29.120 43.710 30.545 43.745 ;
        RECT 44.060 43.710 53.955 43.745 ;
        RECT 44.060 43.705 53.880 43.710 ;
        RECT 44.105 43.685 53.880 43.705 ;
        RECT 53.275 43.640 53.880 43.685 ;
        RECT 34.140 43.255 35.300 43.275 ;
        RECT 44.620 43.255 54.110 43.275 ;
        RECT 26.410 42.715 54.110 43.255 ;
        RECT 26.410 40.225 26.950 42.715 ;
        RECT 27.555 42.185 33.555 42.355 ;
        RECT 27.325 40.975 27.495 42.015 ;
        RECT 33.615 40.975 33.785 42.015 ;
        RECT 27.555 40.635 33.555 40.805 ;
        RECT 34.140 40.225 35.300 42.715 ;
        RECT 42.475 42.695 54.110 42.715 ;
        RECT 35.835 42.185 41.835 42.355 ;
        RECT 35.605 40.975 35.775 42.015 ;
        RECT 41.895 40.975 42.065 42.015 ;
        RECT 35.835 40.635 41.835 40.805 ;
        RECT 42.475 40.290 44.835 42.695 ;
        RECT 45.485 42.185 47.685 42.355 ;
        RECT 45.255 40.975 45.425 42.015 ;
        RECT 47.745 40.975 47.915 42.015 ;
        RECT 45.485 40.635 47.685 40.805 ;
        RECT 48.270 40.290 49.775 42.695 ;
        RECT 50.345 42.190 52.545 42.360 ;
        RECT 50.115 40.980 50.285 42.020 ;
        RECT 52.605 40.980 52.775 42.020 ;
        RECT 50.345 40.640 52.545 40.810 ;
        RECT 53.185 40.290 54.110 42.695 ;
        RECT 42.475 40.225 54.130 40.290 ;
        RECT 26.410 39.455 54.130 40.225 ;
        RECT 26.410 39.180 43.160 39.455 ;
        RECT 53.185 39.430 54.110 39.455 ;
        RECT 26.410 36.670 26.950 39.180 ;
        RECT 27.555 38.605 33.555 38.775 ;
        RECT 27.325 37.395 27.495 38.435 ;
        RECT 33.615 37.395 33.785 38.435 ;
        RECT 27.555 37.055 33.555 37.225 ;
        RECT 34.140 36.670 35.300 39.180 ;
        RECT 35.835 38.605 41.835 38.775 ;
        RECT 35.605 37.395 35.775 38.435 ;
        RECT 41.895 37.395 42.065 38.435 ;
        RECT 35.835 37.055 41.835 37.225 ;
        RECT 42.475 36.670 43.160 39.180 ;
        RECT 26.410 35.625 43.160 36.670 ;
        RECT 26.410 33.050 26.950 35.625 ;
        RECT 27.555 35.025 33.555 35.195 ;
        RECT 27.325 33.815 27.495 34.855 ;
        RECT 33.615 33.815 33.785 34.855 ;
        RECT 27.555 33.475 33.555 33.645 ;
        RECT 34.140 33.050 35.300 35.625 ;
        RECT 35.835 35.025 41.835 35.195 ;
        RECT 35.605 33.815 35.775 34.855 ;
        RECT 41.895 33.815 42.065 34.855 ;
        RECT 35.835 33.475 41.835 33.645 ;
        RECT 42.475 33.050 43.160 35.625 ;
        RECT 26.410 32.005 43.160 33.050 ;
        RECT 26.410 29.555 26.950 32.005 ;
        RECT 27.555 31.445 33.555 31.615 ;
        RECT 27.325 30.235 27.495 31.275 ;
        RECT 33.615 30.235 33.785 31.275 ;
        RECT 27.555 29.895 33.555 30.065 ;
        RECT 34.140 29.555 35.300 32.005 ;
        RECT 35.835 31.445 41.835 31.615 ;
        RECT 35.605 30.235 35.775 31.275 ;
        RECT 41.895 30.235 42.065 31.275 ;
        RECT 35.835 29.895 41.835 30.065 ;
        RECT 42.475 29.555 43.160 32.005 ;
        RECT 26.410 28.545 43.160 29.555 ;
        RECT 42.475 28.525 43.160 28.545 ;
        RECT 68.460 33.345 70.045 53.945 ;
        RECT 70.485 51.325 70.835 53.485 ;
        RECT 70.485 33.825 70.835 35.985 ;
        RECT 71.315 33.345 71.485 53.945 ;
        RECT 71.965 51.325 72.315 53.485 ;
        RECT 71.965 33.825 72.315 35.985 ;
        RECT 72.795 33.345 72.965 53.945 ;
        RECT 73.445 51.325 73.795 53.485 ;
        RECT 73.445 33.825 73.795 35.985 ;
        RECT 74.275 33.345 74.445 53.945 ;
        RECT 74.925 51.325 75.275 53.485 ;
        RECT 74.925 33.825 75.275 35.985 ;
        RECT 75.755 33.345 75.925 53.945 ;
        RECT 76.405 51.325 76.755 53.485 ;
        RECT 76.405 33.825 76.755 35.985 ;
        RECT 77.235 33.345 77.405 53.945 ;
        RECT 77.885 51.325 78.235 53.485 ;
        RECT 77.885 33.825 78.235 35.985 ;
        RECT 78.715 33.345 78.885 53.945 ;
        RECT 79.365 51.325 79.715 53.485 ;
        RECT 79.365 33.825 79.715 35.985 ;
        RECT 80.195 33.345 80.365 53.945 ;
        RECT 80.845 51.325 81.195 53.485 ;
        RECT 81.650 49.365 102.225 53.945 ;
        RECT 81.590 49.150 102.225 49.365 ;
        RECT 81.590 37.665 82.720 49.150 ;
        RECT 83.275 48.630 83.775 48.800 ;
        RECT 84.065 48.630 84.565 48.800 ;
        RECT 84.855 48.630 85.355 48.800 ;
        RECT 85.645 48.630 86.145 48.800 ;
        RECT 86.435 48.630 86.935 48.800 ;
        RECT 87.225 48.630 87.725 48.800 ;
        RECT 88.015 48.630 88.515 48.800 ;
        RECT 88.805 48.630 89.305 48.800 ;
        RECT 89.595 48.630 90.095 48.800 ;
        RECT 90.385 48.630 90.885 48.800 ;
        RECT 91.175 48.630 91.675 48.800 ;
        RECT 91.965 48.630 92.465 48.800 ;
        RECT 92.755 48.630 93.255 48.800 ;
        RECT 93.545 48.630 94.045 48.800 ;
        RECT 94.335 48.630 94.835 48.800 ;
        RECT 95.125 48.630 95.625 48.800 ;
        RECT 95.915 48.630 96.415 48.800 ;
        RECT 96.705 48.630 97.205 48.800 ;
        RECT 97.495 48.630 97.995 48.800 ;
        RECT 98.285 48.630 98.785 48.800 ;
        RECT 99.075 48.630 99.575 48.800 ;
        RECT 99.865 48.630 100.365 48.800 ;
        RECT 83.045 38.420 83.215 48.460 ;
        RECT 83.835 38.420 84.005 48.460 ;
        RECT 84.625 38.420 84.795 48.460 ;
        RECT 85.415 38.420 85.585 48.460 ;
        RECT 86.205 38.420 86.375 48.460 ;
        RECT 86.995 38.420 87.165 48.460 ;
        RECT 87.785 38.420 87.955 48.460 ;
        RECT 88.575 38.420 88.745 48.460 ;
        RECT 89.365 38.420 89.535 48.460 ;
        RECT 90.155 38.420 90.325 48.460 ;
        RECT 90.945 38.420 91.115 48.460 ;
        RECT 91.735 38.420 91.905 48.460 ;
        RECT 92.525 38.420 92.695 48.460 ;
        RECT 93.315 38.420 93.485 48.460 ;
        RECT 94.105 38.420 94.275 48.460 ;
        RECT 94.895 38.420 95.065 48.460 ;
        RECT 95.685 38.420 95.855 48.460 ;
        RECT 96.475 38.420 96.645 48.460 ;
        RECT 97.265 38.420 97.435 48.460 ;
        RECT 98.055 38.420 98.225 48.460 ;
        RECT 98.845 38.420 99.015 48.460 ;
        RECT 99.635 38.420 99.805 48.460 ;
        RECT 100.425 38.420 100.595 48.460 ;
        RECT 83.275 38.080 83.775 38.250 ;
        RECT 84.065 38.080 84.565 38.250 ;
        RECT 84.855 38.080 85.355 38.250 ;
        RECT 85.645 38.080 86.145 38.250 ;
        RECT 86.435 38.080 86.935 38.250 ;
        RECT 87.225 38.080 87.725 38.250 ;
        RECT 88.015 38.080 88.515 38.250 ;
        RECT 88.805 38.080 89.305 38.250 ;
        RECT 89.595 38.080 90.095 38.250 ;
        RECT 90.385 38.080 90.885 38.250 ;
        RECT 91.175 38.080 91.675 38.250 ;
        RECT 91.965 38.080 92.465 38.250 ;
        RECT 92.755 38.080 93.255 38.250 ;
        RECT 93.545 38.080 94.045 38.250 ;
        RECT 94.335 38.080 94.835 38.250 ;
        RECT 95.125 38.080 95.625 38.250 ;
        RECT 95.915 38.080 96.415 38.250 ;
        RECT 96.705 38.080 97.205 38.250 ;
        RECT 97.495 38.080 97.995 38.250 ;
        RECT 98.285 38.080 98.785 38.250 ;
        RECT 99.075 38.080 99.575 38.250 ;
        RECT 99.865 38.080 100.365 38.250 ;
        RECT 100.985 37.665 102.225 49.150 ;
        RECT 81.590 36.320 102.225 37.665 ;
        RECT 80.845 33.825 81.195 35.985 ;
        RECT 81.590 33.345 82.720 36.320 ;
        RECT 83.385 35.715 84.425 35.885 ;
        RECT 68.460 33.175 82.720 33.345 ;
        RECT 68.460 12.700 70.045 33.175 ;
        RECT 70.485 30.535 70.835 32.695 ;
        RECT 70.485 13.035 70.835 15.195 ;
        RECT 71.315 12.700 71.485 33.175 ;
        RECT 71.965 30.535 72.315 32.695 ;
        RECT 71.965 13.035 72.315 15.195 ;
        RECT 72.795 12.700 72.965 33.175 ;
        RECT 73.445 30.535 73.795 32.695 ;
        RECT 73.445 13.035 73.795 15.195 ;
        RECT 74.275 12.700 74.445 33.175 ;
        RECT 74.925 30.535 75.275 32.695 ;
        RECT 74.925 13.035 75.275 15.195 ;
        RECT 75.755 12.700 75.925 33.175 ;
        RECT 76.405 30.535 76.755 32.695 ;
        RECT 76.405 13.035 76.755 15.195 ;
        RECT 77.235 12.700 77.405 33.175 ;
        RECT 77.885 30.535 78.235 32.695 ;
        RECT 77.885 13.035 78.235 15.195 ;
        RECT 78.715 12.700 78.885 33.175 ;
        RECT 79.365 30.535 79.715 32.695 ;
        RECT 79.365 13.035 79.715 15.195 ;
        RECT 80.195 12.700 80.365 33.175 ;
        RECT 80.845 30.535 81.195 32.695 ;
        RECT 81.590 24.925 82.720 33.175 ;
        RECT 83.045 25.655 83.215 35.655 ;
        RECT 84.595 25.655 84.765 35.655 ;
        RECT 83.385 25.425 84.425 25.595 ;
        RECT 85.285 24.925 85.455 36.320 ;
        RECT 86.315 35.715 87.355 35.885 ;
        RECT 85.975 25.655 86.145 35.655 ;
        RECT 87.525 25.655 87.695 35.655 ;
        RECT 86.315 25.425 87.355 25.595 ;
        RECT 88.215 24.925 88.385 36.320 ;
        RECT 89.245 35.715 90.285 35.885 ;
        RECT 88.905 25.655 89.075 35.655 ;
        RECT 90.455 25.655 90.625 35.655 ;
        RECT 91.145 31.650 102.225 36.320 ;
        RECT 89.245 25.425 90.285 25.595 ;
        RECT 91.145 24.925 93.105 31.650 ;
        RECT 93.570 29.035 93.920 31.195 ;
        RECT 81.590 24.755 93.105 24.925 ;
        RECT 81.590 24.245 82.720 24.755 ;
        RECT 91.180 24.245 93.105 24.755 ;
        RECT 81.590 24.075 93.105 24.245 ;
        RECT 80.845 13.035 81.195 15.195 ;
        RECT 81.590 12.700 82.720 24.075 ;
        RECT 83.385 23.405 84.425 23.575 ;
        RECT 83.045 13.345 83.215 23.345 ;
        RECT 84.595 13.345 84.765 23.345 ;
        RECT 83.385 13.115 84.425 13.285 ;
        RECT 85.285 12.700 85.455 24.075 ;
        RECT 86.315 23.405 87.355 23.575 ;
        RECT 85.975 13.345 86.145 23.345 ;
        RECT 87.525 13.345 87.695 23.345 ;
        RECT 86.315 13.115 87.355 13.285 ;
        RECT 88.215 12.700 88.385 24.075 ;
        RECT 89.245 23.405 90.285 23.575 ;
        RECT 88.905 13.345 89.075 23.345 ;
        RECT 90.455 13.345 90.625 23.345 ;
        RECT 89.245 13.115 90.285 13.285 ;
        RECT 91.145 12.700 93.105 24.075 ;
        RECT 93.570 13.035 93.920 15.195 ;
        RECT 94.400 12.700 94.570 31.650 ;
        RECT 95.050 29.035 95.400 31.195 ;
        RECT 95.050 13.035 95.400 15.195 ;
        RECT 95.880 12.700 96.050 31.650 ;
        RECT 96.530 29.035 96.880 31.195 ;
        RECT 96.530 13.035 96.880 15.195 ;
        RECT 97.360 12.700 97.530 31.650 ;
        RECT 98.010 29.035 98.360 31.195 ;
        RECT 98.010 13.035 98.360 15.195 ;
        RECT 98.840 12.700 102.225 31.650 ;
        RECT 68.460 11.055 102.225 12.700 ;
        RECT 105.930 39.940 120.710 40.895 ;
        RECT 105.930 29.855 107.925 39.940 ;
        RECT 108.665 39.555 118.705 39.725 ;
        RECT 108.325 30.495 108.495 39.495 ;
        RECT 118.875 30.495 119.045 39.495 ;
        RECT 108.665 30.265 118.705 30.435 ;
        RECT 119.425 29.855 120.710 39.940 ;
        RECT 105.930 28.940 120.710 29.855 ;
        RECT 105.930 18.625 107.925 28.940 ;
        RECT 108.665 28.305 118.705 28.475 ;
        RECT 108.325 19.245 108.495 28.245 ;
        RECT 118.875 19.245 119.045 28.245 ;
        RECT 119.425 21.810 120.710 28.940 ;
        RECT 121.605 40.170 134.335 40.895 ;
        RECT 121.605 37.835 123.445 40.170 ;
        RECT 124.135 39.555 128.175 39.725 ;
        RECT 123.750 38.495 123.920 39.495 ;
        RECT 128.390 38.495 128.560 39.495 ;
        RECT 124.135 38.265 128.175 38.435 ;
        RECT 129.005 37.835 134.335 40.170 ;
        RECT 121.605 36.585 134.335 37.835 ;
        RECT 121.605 25.405 123.445 36.585 ;
        RECT 124.135 36.025 132.675 36.195 ;
        RECT 123.750 34.965 123.920 35.965 ;
        RECT 132.890 34.965 133.060 35.965 ;
        RECT 124.135 34.735 132.675 34.905 ;
        RECT 123.750 33.675 123.920 34.675 ;
        RECT 132.890 33.675 133.060 34.675 ;
        RECT 124.135 33.445 132.675 33.615 ;
        RECT 123.750 32.385 123.920 33.385 ;
        RECT 132.890 32.385 133.060 33.385 ;
        RECT 124.135 32.155 132.675 32.325 ;
        RECT 123.750 31.095 123.920 32.095 ;
        RECT 132.890 31.095 133.060 32.095 ;
        RECT 124.135 30.865 132.675 31.035 ;
        RECT 123.750 29.805 123.920 30.805 ;
        RECT 132.890 29.805 133.060 30.805 ;
        RECT 124.135 29.575 132.675 29.745 ;
        RECT 123.750 28.515 123.920 29.515 ;
        RECT 132.890 28.515 133.060 29.515 ;
        RECT 124.135 28.285 132.675 28.455 ;
        RECT 123.750 27.225 123.920 28.225 ;
        RECT 132.890 27.225 133.060 28.225 ;
        RECT 124.135 26.995 132.675 27.165 ;
        RECT 123.750 25.935 123.920 26.935 ;
        RECT 132.890 25.935 133.060 26.935 ;
        RECT 124.135 25.705 132.675 25.875 ;
        RECT 133.345 25.405 134.335 36.585 ;
        RECT 121.605 22.245 134.335 25.405 ;
        RECT 119.425 19.685 134.590 21.810 ;
        RECT 108.665 19.015 118.705 19.185 ;
        RECT 119.425 18.625 122.640 19.685 ;
        RECT 123.310 19.015 133.350 19.185 ;
        RECT 105.930 15.415 122.640 18.625 ;
        RECT 105.930 9.025 106.810 15.415 ;
        RECT 107.460 14.825 108.460 14.995 ;
        RECT 108.750 14.825 109.750 14.995 ;
        RECT 110.040 14.825 111.040 14.995 ;
        RECT 111.330 14.825 112.330 14.995 ;
        RECT 112.620 14.825 113.620 14.995 ;
        RECT 113.910 14.825 114.910 14.995 ;
        RECT 115.200 14.825 116.200 14.995 ;
        RECT 116.490 14.825 117.490 14.995 ;
        RECT 117.780 14.825 118.780 14.995 ;
        RECT 119.070 14.825 120.070 14.995 ;
        RECT 107.230 9.615 107.400 14.655 ;
        RECT 108.520 9.615 108.690 14.655 ;
        RECT 109.810 9.615 109.980 14.655 ;
        RECT 111.100 9.615 111.270 14.655 ;
        RECT 112.390 9.615 112.560 14.655 ;
        RECT 113.680 9.615 113.850 14.655 ;
        RECT 114.970 9.615 115.140 14.655 ;
        RECT 116.260 9.615 116.430 14.655 ;
        RECT 117.550 9.615 117.720 14.655 ;
        RECT 118.840 9.615 119.010 14.655 ;
        RECT 120.130 9.615 120.300 14.655 ;
        RECT 107.460 9.275 108.460 9.445 ;
        RECT 108.750 9.275 109.750 9.445 ;
        RECT 110.040 9.275 111.040 9.445 ;
        RECT 111.330 9.275 112.330 9.445 ;
        RECT 112.620 9.275 113.620 9.445 ;
        RECT 113.910 9.275 114.910 9.445 ;
        RECT 115.200 9.275 116.200 9.445 ;
        RECT 116.490 9.275 117.490 9.445 ;
        RECT 117.780 9.275 118.780 9.445 ;
        RECT 119.070 9.275 120.070 9.445 ;
        RECT 120.750 9.435 122.640 15.415 ;
        RECT 122.970 9.955 123.140 18.955 ;
        RECT 133.520 9.955 133.690 18.955 ;
        RECT 123.310 9.725 133.350 9.895 ;
        RECT 134.125 9.435 134.590 19.685 ;
        RECT 120.750 9.025 134.590 9.435 ;
        RECT 105.930 8.145 134.590 9.025 ;
      LAYER met1 ;
        RECT 12.125 212.920 13.435 212.945 ;
        RECT 12.125 212.890 29.205 212.920 ;
        RECT 12.115 211.705 29.205 212.890 ;
        RECT 12.115 151.255 13.490 211.705 ;
        RECT 13.980 210.835 15.710 211.160 ;
        RECT 13.980 209.055 14.230 210.835 ;
        RECT 15.460 209.055 15.710 210.835 ;
        RECT 16.940 210.835 18.670 211.160 ;
        RECT 16.940 209.055 17.190 210.835 ;
        RECT 18.420 209.055 18.670 210.835 ;
        RECT 19.900 210.835 21.630 211.160 ;
        RECT 19.900 209.055 20.150 210.835 ;
        RECT 21.380 209.055 21.630 210.835 ;
        RECT 22.860 210.835 24.590 211.160 ;
        RECT 22.860 209.055 23.110 210.835 ;
        RECT 24.340 209.055 24.590 210.835 ;
        RECT 25.820 210.835 27.550 211.160 ;
        RECT 25.820 209.055 26.070 210.835 ;
        RECT 27.300 209.055 27.550 210.835 ;
        RECT 13.980 178.765 14.230 184.165 ;
        RECT 15.460 178.765 15.710 184.165 ;
        RECT 16.940 178.765 17.190 184.165 ;
        RECT 18.420 178.765 18.670 184.165 ;
        RECT 19.900 178.765 20.150 184.165 ;
        RECT 21.380 178.765 21.630 184.165 ;
        RECT 22.860 178.765 23.110 184.165 ;
        RECT 24.340 178.765 24.590 184.165 ;
        RECT 25.820 178.765 26.070 184.165 ;
        RECT 27.300 178.765 27.550 184.165 ;
        RECT 27.965 155.000 29.125 211.705 ;
        RECT 30.100 155.560 54.475 156.545 ;
        RECT 13.980 153.830 14.230 153.875 ;
        RECT 13.870 151.830 14.330 153.830 ;
        RECT 15.460 152.095 15.710 153.875 ;
        RECT 16.940 152.095 17.190 153.875 ;
        RECT 13.980 151.770 14.230 151.830 ;
        RECT 15.460 151.770 17.190 152.095 ;
        RECT 18.420 152.095 18.670 153.875 ;
        RECT 19.900 152.095 20.150 153.875 ;
        RECT 18.420 151.770 20.150 152.095 ;
        RECT 21.380 152.095 21.630 153.875 ;
        RECT 22.860 152.095 23.110 153.875 ;
        RECT 21.380 151.770 23.110 152.095 ;
        RECT 24.340 152.095 24.590 153.875 ;
        RECT 25.820 152.095 26.070 153.875 ;
        RECT 27.300 153.815 27.550 153.875 ;
        RECT 24.340 151.770 26.070 152.095 ;
        RECT 27.245 151.830 27.605 153.815 ;
        RECT 27.300 151.770 27.550 151.830 ;
        RECT 28.035 151.255 29.105 155.000 ;
        RECT 30.110 152.710 30.745 155.560 ;
        RECT 31.415 154.795 41.375 155.025 ;
        RECT 43.045 154.795 53.005 155.025 ;
        RECT 31.135 154.150 31.365 154.590 ;
        RECT 31.070 153.650 31.430 154.150 ;
        RECT 41.425 153.920 41.655 154.590 ;
        RECT 42.765 153.920 42.995 154.590 ;
        RECT 53.055 154.530 53.285 154.590 ;
        RECT 52.960 154.030 53.380 154.530 ;
        RECT 31.135 153.590 31.365 153.650 ;
        RECT 41.425 153.590 42.995 153.920 ;
        RECT 53.055 153.590 53.285 154.030 ;
        RECT 31.425 153.385 32.790 153.395 ;
        RECT 51.095 153.385 52.995 153.430 ;
        RECT 31.415 153.155 53.005 153.385 ;
        RECT 31.425 153.110 32.790 153.155 ;
        RECT 51.095 153.065 52.995 153.155 ;
        RECT 53.745 152.710 54.420 155.560 ;
        RECT 30.095 151.725 54.470 152.710 ;
        RECT 12.115 151.250 29.135 151.255 ;
        RECT 12.095 150.315 29.135 151.250 ;
        RECT 12.125 150.260 29.135 150.315 ;
        RECT 12.125 150.255 13.435 150.260 ;
        RECT 36.790 140.920 88.970 141.775 ;
        RECT 36.790 140.515 37.480 140.920 ;
        RECT 66.995 140.840 88.970 140.920 ;
        RECT 66.995 140.515 88.020 140.840 ;
        RECT 36.790 140.265 40.065 140.515 ;
        RECT 49.455 140.265 88.020 140.515 ;
        RECT 36.790 139.925 37.480 140.265 ;
        RECT 35.520 139.915 37.480 139.925 ;
        RECT 31.130 137.910 37.480 139.915 ;
        RECT 66.995 140.220 88.020 140.265 ;
        RECT 64.255 139.035 66.340 139.040 ;
        RECT 36.790 124.285 37.480 137.910 ;
        RECT 37.960 138.785 40.065 139.035 ;
        RECT 49.455 138.785 54.855 139.035 ;
        RECT 64.245 138.785 66.350 139.035 ;
        RECT 37.960 137.555 38.370 138.785 ;
        RECT 64.255 138.780 66.340 138.785 ;
        RECT 37.960 137.305 40.065 137.555 ;
        RECT 49.455 137.305 54.855 137.555 ;
        RECT 64.245 137.305 66.350 137.555 ;
        RECT 65.940 136.075 66.350 137.305 ;
        RECT 37.960 135.825 40.065 136.075 ;
        RECT 49.455 135.825 54.855 136.075 ;
        RECT 64.245 135.825 66.350 136.075 ;
        RECT 66.995 135.920 69.250 140.220 ;
        RECT 69.930 139.090 72.980 139.615 ;
        RECT 73.635 139.095 75.965 140.220 ;
        RECT 69.880 138.750 72.980 139.090 ;
        RECT 76.650 138.750 79.700 139.615 ;
        RECT 80.360 139.040 82.690 140.220 ;
        RECT 69.880 138.720 79.700 138.750 ;
        RECT 83.370 138.720 86.420 139.615 ;
        RECT 69.880 137.350 86.420 138.720 ;
        RECT 69.880 136.720 72.980 137.350 ;
        RECT 76.650 137.320 86.420 137.350 ;
        RECT 69.930 136.565 72.980 136.720 ;
        RECT 37.960 134.595 38.370 135.825 ;
        RECT 37.960 134.345 40.065 134.595 ;
        RECT 49.455 134.345 54.855 134.595 ;
        RECT 64.245 134.345 66.350 134.595 ;
        RECT 65.940 133.115 66.350 134.345 ;
        RECT 37.960 132.865 40.065 133.115 ;
        RECT 49.455 132.865 54.855 133.115 ;
        RECT 64.245 132.865 66.350 133.115 ;
        RECT 66.995 134.255 70.440 135.920 ;
        RECT 37.960 131.635 38.370 132.865 ;
        RECT 37.960 131.385 40.065 131.635 ;
        RECT 49.455 131.385 54.855 131.635 ;
        RECT 64.245 131.385 66.350 131.635 ;
        RECT 65.940 130.155 66.350 131.385 ;
        RECT 37.960 129.905 40.065 130.155 ;
        RECT 49.455 129.905 54.855 130.155 ;
        RECT 64.245 129.905 66.350 130.155 ;
        RECT 37.960 128.675 38.370 129.905 ;
        RECT 66.995 129.190 69.250 134.255 ;
        RECT 70.715 132.895 72.260 136.565 ;
        RECT 73.780 135.905 75.920 136.920 ;
        RECT 76.650 136.565 79.700 137.320 ;
        RECT 80.430 135.905 82.570 136.920 ;
        RECT 83.370 136.565 86.420 137.320 ;
        RECT 72.690 134.355 83.880 135.905 ;
        RECT 69.930 129.845 72.980 132.895 ;
        RECT 37.960 128.425 40.065 128.675 ;
        RECT 49.455 128.425 54.855 128.675 ;
        RECT 64.245 128.425 66.350 128.675 ;
        RECT 65.940 127.195 66.350 128.425 ;
        RECT 37.960 126.945 40.065 127.195 ;
        RECT 49.455 126.945 54.855 127.195 ;
        RECT 64.245 126.945 66.350 127.195 ;
        RECT 66.995 127.525 70.440 129.190 ;
        RECT 37.960 125.715 38.370 126.945 ;
        RECT 64.740 125.715 66.340 125.720 ;
        RECT 37.960 125.465 40.065 125.715 ;
        RECT 49.455 125.465 54.855 125.715 ;
        RECT 64.245 125.465 66.350 125.715 ;
        RECT 64.740 125.460 66.340 125.465 ;
        RECT 36.790 124.235 38.060 124.285 ;
        RECT 66.995 124.240 69.250 127.525 ;
        RECT 70.700 126.175 72.245 129.845 ;
        RECT 73.780 129.160 75.920 134.355 ;
        RECT 76.650 129.845 79.700 132.895 ;
        RECT 80.430 129.160 82.570 134.355 ;
        RECT 84.195 132.895 85.740 136.565 ;
        RECT 87.090 135.955 88.020 140.220 ;
        RECT 85.945 134.290 88.020 135.955 ;
        RECT 83.370 129.845 86.420 132.895 ;
        RECT 72.845 127.570 83.825 129.160 ;
        RECT 66.280 124.235 69.250 124.240 ;
        RECT 36.790 123.985 69.250 124.235 ;
        RECT 36.790 123.935 38.060 123.985 ;
        RECT 28.680 123.135 29.935 123.165 ;
        RECT 36.790 123.135 37.480 123.935 ;
        RECT 28.680 123.105 37.480 123.135 ;
        RECT 28.660 123.100 37.480 123.105 ;
        RECT 66.995 123.100 69.250 123.985 ;
        RECT 69.930 125.250 72.980 126.175 ;
        RECT 73.780 125.465 75.920 127.570 ;
        RECT 76.650 125.250 79.700 126.175 ;
        RECT 80.430 125.465 82.570 127.570 ;
        RECT 84.220 126.175 85.765 129.845 ;
        RECT 87.090 129.285 88.020 134.290 ;
        RECT 86.020 127.445 88.020 129.285 ;
        RECT 69.930 125.235 79.700 125.250 ;
        RECT 83.370 125.235 86.420 126.175 ;
        RECT 69.930 123.850 86.420 125.235 ;
        RECT 69.930 123.125 72.980 123.850 ;
        RECT 76.650 123.835 86.420 123.850 ;
        RECT 28.660 122.510 69.250 123.100 ;
        RECT 73.655 122.510 75.985 123.610 ;
        RECT 76.650 123.125 79.700 123.835 ;
        RECT 80.380 122.510 82.710 123.590 ;
        RECT 83.370 123.125 86.420 123.835 ;
        RECT 87.090 122.510 88.020 127.445 ;
        RECT 28.660 121.965 88.020 122.510 ;
        RECT 28.660 120.960 88.050 121.965 ;
        RECT 28.660 99.800 29.955 120.960 ;
        RECT 30.760 120.510 31.260 120.540 ;
        RECT 30.740 120.340 31.280 120.510 ;
        RECT 30.760 120.310 31.260 120.340 ;
        RECT 30.370 118.870 30.600 120.285 ;
        RECT 30.850 120.250 31.250 120.310 ;
        RECT 31.420 119.805 31.650 120.280 ;
        RECT 31.350 118.870 31.710 119.805 ;
        RECT 30.370 114.805 31.710 118.870 ;
        RECT 30.370 101.660 31.650 114.805 ;
        RECT 30.370 100.220 30.600 101.660 ;
        RECT 30.760 100.220 31.260 100.250 ;
        RECT 31.420 100.220 31.650 101.660 ;
        RECT 30.370 100.050 31.650 100.220 ;
        RECT 30.760 100.020 31.260 100.050 ;
        RECT 30.850 99.990 31.250 100.020 ;
        RECT 32.110 99.800 32.340 120.960 ;
        RECT 33.190 120.310 33.690 120.540 ;
        RECT 32.800 119.805 33.030 120.260 ;
        RECT 33.200 120.250 33.600 120.310 ;
        RECT 33.850 119.805 34.080 120.260 ;
        RECT 32.740 118.870 33.100 119.805 ;
        RECT 33.790 118.870 34.150 119.805 ;
        RECT 32.740 114.805 34.150 118.870 ;
        RECT 32.800 101.660 34.080 114.805 ;
        RECT 32.800 100.300 33.030 101.660 ;
        RECT 33.850 100.300 34.080 101.660 ;
        RECT 33.190 100.020 33.690 100.250 ;
        RECT 33.280 99.960 33.680 100.020 ;
        RECT 34.540 99.800 34.770 120.960 ;
        RECT 35.710 120.540 36.110 120.600 ;
        RECT 35.620 120.310 36.120 120.540 ;
        RECT 35.230 119.815 35.460 120.260 ;
        RECT 35.180 118.870 35.540 119.815 ;
        RECT 36.280 118.870 36.510 120.260 ;
        RECT 35.180 114.815 36.510 118.870 ;
        RECT 35.230 101.660 36.510 114.815 ;
        RECT 35.230 100.300 35.460 101.660 ;
        RECT 36.280 100.300 36.510 101.660 ;
        RECT 35.620 100.020 36.120 100.250 ;
        RECT 35.630 99.960 36.030 100.020 ;
        RECT 36.970 99.800 37.200 120.960 ;
        RECT 38.140 120.540 38.540 120.600 ;
        RECT 38.050 120.510 38.550 120.540 ;
        RECT 38.050 120.340 38.570 120.510 ;
        RECT 38.050 120.310 38.550 120.340 ;
        RECT 37.660 118.915 37.890 120.280 ;
        RECT 38.710 119.830 38.940 120.290 ;
        RECT 38.635 118.915 38.995 119.830 ;
        RECT 37.660 114.830 38.995 118.915 ;
        RECT 37.660 101.685 38.940 114.830 ;
        RECT 37.660 100.220 37.890 101.685 ;
        RECT 38.050 100.220 38.550 100.250 ;
        RECT 38.710 100.220 38.940 101.685 ;
        RECT 37.660 100.050 38.940 100.220 ;
        RECT 38.050 100.045 38.940 100.050 ;
        RECT 38.050 100.020 38.550 100.045 ;
        RECT 38.060 99.960 38.460 100.020 ;
        RECT 39.400 99.800 39.630 120.960 ;
        RECT 40.490 120.540 40.890 120.600 ;
        RECT 40.480 120.310 40.980 120.540 ;
        RECT 40.090 119.830 40.320 120.260 ;
        RECT 40.030 118.915 40.390 119.830 ;
        RECT 41.140 119.820 41.370 120.260 ;
        RECT 41.075 118.915 41.435 119.820 ;
        RECT 40.030 114.830 41.435 118.915 ;
        RECT 40.090 114.820 41.435 114.830 ;
        RECT 40.090 101.685 41.370 114.820 ;
        RECT 40.090 100.300 40.320 101.685 ;
        RECT 41.140 100.300 41.370 101.685 ;
        RECT 40.480 100.020 40.980 100.250 ;
        RECT 40.570 99.960 40.970 100.020 ;
        RECT 41.830 99.800 42.060 120.960 ;
        RECT 43.000 120.540 43.400 120.600 ;
        RECT 42.910 120.310 43.410 120.540 ;
        RECT 42.520 119.820 42.750 120.260 ;
        RECT 42.450 118.930 42.810 119.820 ;
        RECT 43.570 119.815 43.800 120.260 ;
        RECT 43.510 118.930 43.870 119.815 ;
        RECT 42.450 114.820 43.870 118.930 ;
        RECT 42.520 114.815 43.870 114.820 ;
        RECT 42.520 101.700 43.800 114.815 ;
        RECT 42.520 100.300 42.750 101.700 ;
        RECT 43.570 100.300 43.800 101.700 ;
        RECT 42.910 100.020 43.410 100.250 ;
        RECT 42.920 99.960 43.320 100.020 ;
        RECT 44.260 99.800 44.490 120.960 ;
        RECT 45.350 120.540 45.750 120.600 ;
        RECT 45.340 120.310 45.840 120.540 ;
        RECT 44.950 119.815 45.180 120.260 ;
        RECT 46.000 119.815 46.230 120.260 ;
        RECT 44.885 118.930 45.245 119.815 ;
        RECT 45.935 118.930 46.295 119.815 ;
        RECT 44.885 114.815 46.295 118.930 ;
        RECT 44.950 101.700 46.230 114.815 ;
        RECT 44.950 100.300 45.180 101.700 ;
        RECT 46.000 100.300 46.230 101.700 ;
        RECT 45.340 100.020 45.840 100.250 ;
        RECT 45.430 99.960 45.830 100.020 ;
        RECT 46.690 99.800 46.920 120.960 ;
        RECT 47.860 120.540 48.260 120.600 ;
        RECT 47.770 120.310 48.270 120.540 ;
        RECT 47.380 119.815 47.610 120.260 ;
        RECT 48.430 119.815 48.660 120.260 ;
        RECT 47.315 118.930 47.675 119.815 ;
        RECT 48.370 118.930 48.730 119.815 ;
        RECT 47.315 114.815 48.730 118.930 ;
        RECT 47.380 101.700 48.660 114.815 ;
        RECT 47.380 100.300 47.610 101.700 ;
        RECT 48.430 100.300 48.660 101.700 ;
        RECT 47.770 100.020 48.270 100.250 ;
        RECT 47.780 99.960 48.180 100.020 ;
        RECT 49.120 99.800 49.350 120.960 ;
        RECT 50.210 120.540 50.610 120.600 ;
        RECT 50.200 120.310 50.700 120.540 ;
        RECT 49.810 119.815 50.040 120.260 ;
        RECT 50.860 119.815 51.090 120.260 ;
        RECT 49.745 118.930 50.105 119.815 ;
        RECT 50.795 118.930 51.155 119.815 ;
        RECT 49.745 114.815 51.155 118.930 ;
        RECT 49.810 101.700 51.090 114.815 ;
        RECT 49.810 100.300 50.040 101.700 ;
        RECT 50.860 100.300 51.090 101.700 ;
        RECT 50.200 100.020 50.700 100.250 ;
        RECT 50.290 99.960 50.690 100.020 ;
        RECT 51.550 99.800 51.780 120.960 ;
        RECT 52.720 120.540 53.120 120.600 ;
        RECT 52.630 120.310 53.130 120.540 ;
        RECT 52.240 119.815 52.470 120.260 ;
        RECT 52.180 118.945 52.540 119.815 ;
        RECT 53.290 118.945 53.520 120.260 ;
        RECT 52.180 114.815 53.520 118.945 ;
        RECT 52.240 101.715 53.520 114.815 ;
        RECT 52.240 100.300 52.470 101.715 ;
        RECT 53.290 100.300 53.520 101.715 ;
        RECT 53.825 117.610 54.305 120.960 ;
        RECT 77.745 120.275 88.050 120.960 ;
        RECT 99.795 120.275 100.775 120.305 ;
        RECT 77.745 118.885 100.775 120.275 ;
        RECT 79.235 118.255 99.195 118.485 ;
        RECT 78.955 118.035 79.185 118.095 ;
        RECT 53.825 117.580 54.730 117.610 ;
        RECT 53.825 116.790 78.035 117.580 ;
        RECT 78.890 117.035 79.250 118.035 ;
        RECT 53.825 116.760 54.730 116.790 ;
        RECT 53.825 116.755 54.620 116.760 ;
        RECT 53.825 103.980 54.305 116.755 ;
        RECT 55.340 111.810 56.130 116.790 ;
        RECT 56.705 116.255 76.915 116.485 ;
        RECT 56.705 116.095 56.875 116.255 ;
        RECT 56.675 114.155 56.905 116.095 ;
        RECT 56.610 113.155 56.970 114.155 ;
        RECT 56.675 113.095 56.905 113.155 ;
        RECT 56.705 112.935 56.875 113.095 ;
        RECT 65.180 112.935 69.430 116.255 ;
        RECT 76.965 114.155 77.195 116.095 ;
        RECT 76.900 113.155 77.260 114.155 ;
        RECT 76.965 113.095 77.195 113.155 ;
        RECT 78.955 113.095 79.185 117.035 ;
        RECT 87.360 112.935 91.630 118.255 ;
        RECT 99.245 118.035 99.475 118.095 ;
        RECT 99.180 117.035 99.540 118.035 ;
        RECT 99.245 113.095 99.475 117.035 ;
        RECT 56.705 112.705 99.195 112.935 ;
        RECT 75.915 112.390 80.235 112.705 ;
        RECT 55.340 110.830 75.690 111.810 ;
        RECT 55.340 110.800 56.335 110.830 ;
        RECT 53.825 103.950 54.345 103.980 ;
        RECT 55.970 103.950 56.335 110.800 ;
        RECT 75.915 110.440 76.915 112.390 ;
        RECT 79.235 110.440 80.235 112.390 ;
        RECT 99.795 111.965 100.775 118.885 ;
        RECT 80.675 110.700 100.775 111.965 ;
        RECT 75.915 110.125 80.235 110.440 ;
        RECT 56.990 109.895 99.195 110.125 ;
        RECT 56.710 105.795 56.940 109.735 ;
        RECT 56.645 104.795 57.005 105.795 ;
        RECT 56.710 104.735 56.940 104.795 ;
        RECT 65.125 104.575 69.395 109.895 ;
        RECT 78.985 109.735 79.155 109.895 ;
        RECT 77.000 105.795 77.230 109.735 ;
        RECT 78.955 109.675 79.185 109.735 ;
        RECT 77.620 108.840 78.460 108.900 ;
        RECT 77.600 105.975 78.480 108.840 ;
        RECT 78.890 108.675 79.250 109.675 ;
        RECT 78.955 106.735 79.185 108.675 ;
        RECT 78.985 106.575 79.155 106.735 ;
        RECT 87.485 106.575 91.735 109.895 ;
        RECT 99.245 109.675 99.475 109.735 ;
        RECT 99.180 108.675 99.540 109.675 ;
        RECT 99.795 108.760 100.775 110.700 ;
        RECT 99.245 106.735 99.475 108.675 ;
        RECT 78.985 106.345 99.195 106.575 ;
        RECT 99.755 105.975 100.790 108.760 ;
        RECT 76.935 104.795 77.295 105.795 ;
        RECT 77.600 105.550 100.790 105.975 ;
        RECT 77.600 105.375 100.775 105.550 ;
        RECT 77.000 104.735 77.230 104.795 ;
        RECT 56.990 104.345 76.950 104.575 ;
        RECT 53.825 103.945 56.375 103.950 ;
        RECT 77.630 103.945 78.030 105.375 ;
        RECT 99.795 105.345 100.775 105.375 ;
        RECT 53.825 103.450 78.075 103.945 ;
        RECT 52.630 100.020 53.130 100.250 ;
        RECT 52.640 99.960 53.040 100.020 ;
        RECT 53.825 99.800 54.345 103.450 ;
        RECT 55.970 103.420 56.335 103.450 ;
        RECT 77.630 103.435 78.030 103.450 ;
        RECT 28.650 98.625 54.345 99.800 ;
        RECT 30.650 96.200 100.530 96.890 ;
        RECT 30.650 84.405 31.290 96.200 ;
        RECT 46.700 95.690 51.800 95.715 ;
        RECT 32.040 95.460 52.020 95.690 ;
        RECT 33.715 95.435 51.800 95.460 ;
        RECT 31.760 95.195 31.990 95.255 ;
        RECT 31.695 93.815 32.055 95.195 ;
        RECT 31.760 93.755 31.990 93.815 ;
        RECT 33.715 93.550 50.595 95.435 ;
        RECT 52.050 95.195 52.280 95.255 ;
        RECT 51.985 93.815 52.345 95.195 ;
        RECT 52.050 93.755 52.280 93.815 ;
        RECT 32.040 93.320 52.000 93.550 ;
        RECT 32.570 93.010 51.825 93.320 ;
        RECT 32.040 92.780 52.000 93.010 ;
        RECT 31.760 92.515 31.990 92.575 ;
        RECT 31.695 91.135 32.055 92.515 ;
        RECT 31.760 91.075 31.990 91.135 ;
        RECT 33.690 90.870 50.540 92.780 ;
        RECT 52.050 92.515 52.280 92.575 ;
        RECT 51.985 91.135 52.345 92.515 ;
        RECT 52.050 91.075 52.280 91.135 ;
        RECT 32.040 90.640 52.000 90.870 ;
        RECT 49.560 88.690 51.455 90.640 ;
        RECT 32.040 88.460 52.000 88.690 ;
        RECT 31.760 88.195 31.990 88.255 ;
        RECT 31.660 87.195 32.080 88.195 ;
        RECT 31.760 85.255 31.990 87.195 ;
        RECT 33.330 85.050 50.195 88.460 ;
        RECT 52.050 88.195 52.280 88.255 ;
        RECT 51.985 85.315 52.345 88.195 ;
        RECT 52.050 85.255 52.280 85.315 ;
        RECT 32.040 84.820 52.020 85.050 ;
        RECT 39.905 84.405 41.245 84.430 ;
        RECT 52.840 84.405 56.725 96.200 ;
        RECT 57.480 95.690 62.580 95.715 ;
        RECT 57.460 95.460 99.350 95.690 ;
        RECT 57.480 95.435 62.580 95.460 ;
        RECT 57.200 88.315 57.430 95.255 ;
        RECT 57.105 85.315 57.525 88.315 ;
        RECT 57.200 85.255 57.430 85.315 ;
        RECT 65.265 85.050 71.160 95.460 ;
        RECT 77.490 94.645 77.720 95.255 ;
        RECT 78.830 94.645 79.060 95.255 ;
        RECT 77.490 87.815 79.060 94.645 ;
        RECT 77.425 85.775 79.125 87.815 ;
        RECT 77.425 85.315 77.785 85.775 ;
        RECT 78.765 85.315 79.125 85.775 ;
        RECT 77.490 85.255 77.720 85.315 ;
        RECT 78.830 85.255 79.060 85.315 ;
        RECT 86.525 85.050 92.420 95.460 ;
        RECT 99.120 95.195 99.350 95.460 ;
        RECT 99.025 92.195 99.445 95.195 ;
        RECT 99.825 94.990 100.530 96.200 ;
        RECT 99.825 94.265 109.215 94.990 ;
        RECT 99.120 85.255 99.350 92.195 ;
        RECT 99.150 85.050 99.320 85.255 ;
        RECT 57.460 84.820 99.320 85.050 ;
        RECT 30.620 83.675 56.725 84.405 ;
        RECT 30.675 83.665 31.290 83.675 ;
        RECT 40.250 75.175 56.725 83.675 ;
        RECT 57.525 83.670 77.070 84.820 ;
        RECT 79.470 83.670 99.015 84.820 ;
        RECT 57.200 83.440 99.070 83.670 ;
        RECT 57.200 83.175 57.430 83.440 ;
        RECT 57.105 80.175 57.525 83.175 ;
        RECT 40.250 73.945 41.245 75.175 ;
        RECT 42.050 74.670 47.150 74.685 ;
        RECT 42.050 74.440 52.000 74.670 ;
        RECT 42.050 74.425 51.020 74.440 ;
        RECT 40.220 72.350 41.280 73.945 ;
        RECT 41.810 73.930 42.040 74.235 ;
        RECT 41.695 73.295 42.055 73.930 ;
        RECT 41.810 73.235 42.040 73.295 ;
        RECT 43.415 73.030 51.020 74.425 ;
        RECT 52.050 74.175 52.280 74.235 ;
        RECT 51.985 73.295 52.345 74.175 ;
        RECT 52.050 73.235 52.280 73.295 ;
        RECT 42.090 72.800 52.000 73.030 ;
        RECT 52.840 72.350 56.725 75.175 ;
        RECT 57.200 73.235 57.430 80.175 ;
        RECT 57.230 73.030 57.430 73.235 ;
        RECT 65.095 73.030 70.990 83.440 ;
        RECT 77.490 83.175 77.720 83.235 ;
        RECT 78.830 83.175 79.060 83.235 ;
        RECT 77.425 82.655 77.785 83.175 ;
        RECT 78.765 82.655 79.125 83.175 ;
        RECT 77.425 80.675 79.125 82.655 ;
        RECT 77.490 74.250 79.060 80.675 ;
        RECT 77.425 73.725 79.125 74.250 ;
        RECT 77.425 73.295 77.785 73.725 ;
        RECT 78.765 73.295 79.125 73.725 ;
        RECT 77.490 73.235 77.720 73.295 ;
        RECT 78.830 73.235 79.060 73.295 ;
        RECT 86.610 73.030 92.505 83.440 ;
        RECT 99.120 76.295 99.350 83.235 ;
        RECT 99.025 73.890 99.445 76.295 ;
        RECT 99.120 73.235 99.350 73.890 ;
        RECT 57.230 72.800 99.070 73.030 ;
        RECT 99.825 72.350 103.620 94.265 ;
        RECT 104.505 93.870 104.985 93.900 ;
        RECT 104.495 93.640 104.995 93.870 ;
        RECT 106.965 93.660 107.565 93.980 ;
        RECT 107.015 93.640 107.515 93.660 ;
        RECT 104.060 90.345 104.290 93.590 ;
        RECT 105.200 93.500 105.430 93.590 ;
        RECT 105.125 90.345 105.505 93.500 ;
        RECT 104.060 88.500 105.505 90.345 ;
        RECT 106.580 90.345 106.810 93.590 ;
        RECT 107.720 93.290 107.950 93.590 ;
        RECT 107.645 90.345 108.025 93.290 ;
        RECT 104.060 77.360 105.430 88.500 ;
        RECT 104.060 73.630 104.290 77.360 ;
        RECT 105.200 73.630 105.430 77.360 ;
        RECT 106.580 88.290 108.025 90.345 ;
        RECT 106.580 77.360 107.950 88.290 ;
        RECT 106.580 73.630 106.810 77.360 ;
        RECT 107.720 73.630 107.950 77.360 ;
        RECT 104.495 73.350 104.995 73.580 ;
        RECT 107.015 73.350 107.515 73.580 ;
        RECT 104.505 73.320 104.985 73.350 ;
        RECT 107.025 73.320 107.505 73.350 ;
        RECT 108.410 72.350 109.215 94.265 ;
        RECT 40.220 69.945 109.215 72.350 ;
        RECT 38.940 62.565 53.950 64.150 ;
        RECT 29.170 59.875 29.945 59.905 ;
        RECT 38.950 59.875 40.025 62.565 ;
        RECT 40.615 61.820 50.625 62.050 ;
        RECT 40.270 60.675 40.630 61.675 ;
        RECT 40.335 60.615 40.565 60.675 ;
        RECT 42.180 60.420 48.925 61.820 ;
        RECT 50.675 61.555 50.905 61.615 ;
        RECT 50.560 60.675 50.920 61.555 ;
        RECT 50.675 60.615 50.905 60.675 ;
        RECT 40.625 60.410 48.925 60.420 ;
        RECT 40.615 60.180 50.625 60.410 ;
        RECT 40.625 60.160 44.270 60.180 ;
        RECT 51.370 59.875 53.945 62.565 ;
        RECT 29.170 59.845 53.945 59.875 ;
        RECT 29.130 58.755 53.945 59.845 ;
        RECT 29.130 55.970 29.965 58.755 ;
        RECT 30.615 58.005 50.575 58.235 ;
        RECT 30.335 57.740 30.565 57.800 ;
        RECT 29.170 54.940 29.945 55.970 ;
        RECT 30.240 55.860 30.630 57.740 ;
        RECT 30.335 55.800 30.565 55.860 ;
        RECT 35.125 55.595 47.370 58.005 ;
        RECT 50.625 57.740 50.855 57.800 ;
        RECT 50.560 55.860 50.920 57.740 ;
        RECT 50.625 55.800 50.855 55.860 ;
        RECT 30.615 55.365 50.575 55.595 ;
        RECT 30.625 55.315 35.725 55.365 ;
        RECT 51.370 54.940 53.945 58.755 ;
        RECT 59.210 55.615 59.865 55.630 ;
        RECT 59.210 55.570 64.555 55.615 ;
        RECT 29.170 54.780 53.945 54.940 ;
        RECT 29.150 54.200 53.945 54.780 ;
        RECT 29.170 54.030 53.945 54.200 ;
        RECT 59.190 55.000 64.555 55.570 ;
        RECT 68.735 55.240 69.395 55.270 ;
        RECT 68.735 55.160 102.145 55.240 ;
        RECT 29.170 53.975 53.930 54.030 ;
        RECT 29.170 53.945 30.355 53.975 ;
        RECT 29.190 44.385 30.355 53.945 ;
        RECT 31.175 53.075 33.535 53.305 ;
        RECT 35.855 53.075 38.215 53.305 ;
        RECT 30.895 52.810 31.125 52.870 ;
        RECT 30.800 51.635 31.220 52.810 ;
        RECT 30.895 50.370 31.125 51.635 ;
        RECT 31.830 50.165 32.790 53.075 ;
        RECT 33.585 50.960 33.815 52.870 ;
        RECT 34.410 50.960 34.975 50.970 ;
        RECT 35.575 50.960 35.805 52.870 ;
        RECT 33.585 50.370 35.805 50.960 ;
        RECT 31.175 49.935 33.535 50.165 ;
        RECT 31.175 49.590 31.675 49.935 ;
        RECT 34.410 49.850 34.975 50.370 ;
        RECT 36.565 50.165 37.525 53.075 ;
        RECT 38.265 51.610 38.495 52.870 ;
        RECT 38.170 50.430 38.590 51.610 ;
        RECT 38.265 50.370 38.495 50.430 ;
        RECT 35.855 49.965 38.215 50.165 ;
        RECT 35.855 49.935 38.245 49.965 ;
        RECT 31.125 49.090 31.725 49.590 ;
        RECT 32.985 48.340 33.585 48.840 ;
        RECT 33.035 48.095 33.535 48.340 ;
        RECT 31.175 47.865 33.535 48.095 ;
        RECT 30.895 46.400 31.125 47.660 ;
        RECT 30.800 45.220 31.220 46.400 ;
        RECT 30.895 45.160 31.125 45.220 ;
        RECT 31.830 44.955 32.790 47.865 ;
        RECT 34.430 47.660 34.930 49.850 ;
        RECT 35.805 49.090 36.405 49.590 ;
        RECT 35.855 48.095 36.355 49.090 ;
        RECT 37.745 48.840 38.245 49.935 ;
        RECT 37.695 48.340 38.295 48.840 ;
        RECT 35.855 47.865 38.215 48.095 ;
        RECT 33.585 47.070 35.805 47.660 ;
        RECT 33.585 45.160 33.815 47.070 ;
        RECT 35.575 45.160 35.805 47.070 ;
        RECT 36.540 44.955 37.500 47.865 ;
        RECT 38.265 47.600 38.495 47.660 ;
        RECT 38.170 46.425 38.590 47.600 ;
        RECT 38.265 45.160 38.495 46.425 ;
        RECT 31.175 44.725 33.535 44.955 ;
        RECT 35.855 44.725 38.215 44.955 ;
        RECT 38.885 44.385 39.760 53.975 ;
        RECT 29.190 43.805 39.860 44.385 ;
        RECT 44.010 44.345 44.800 53.975 ;
        RECT 51.390 53.970 53.930 53.975 ;
        RECT 45.505 53.165 47.865 53.395 ;
        RECT 50.165 53.165 52.775 53.395 ;
        RECT 45.225 51.520 45.455 52.960 ;
        RECT 45.130 50.520 45.550 51.520 ;
        RECT 45.225 50.460 45.455 50.520 ;
        RECT 45.965 50.255 47.220 53.165 ;
        RECT 47.915 52.900 48.145 52.960 ;
        RECT 49.885 52.900 50.115 52.960 ;
        RECT 47.850 51.900 48.210 52.900 ;
        RECT 49.820 51.900 50.180 52.900 ;
        RECT 47.915 50.460 48.145 51.900 ;
        RECT 49.885 50.460 50.115 51.900 ;
        RECT 50.830 50.255 51.870 53.165 ;
        RECT 52.605 52.960 52.775 53.165 ;
        RECT 52.575 52.900 52.805 52.960 ;
        RECT 52.480 51.900 52.900 52.900 ;
        RECT 52.575 50.460 52.805 51.900 ;
        RECT 52.605 50.255 52.775 50.460 ;
        RECT 45.505 50.225 47.865 50.255 ;
        RECT 50.165 50.225 52.775 50.255 ;
        RECT 45.505 50.055 52.775 50.225 ;
        RECT 45.505 50.025 47.865 50.055 ;
        RECT 47.240 47.970 47.865 50.025 ;
        RECT 45.255 47.940 47.865 47.970 ;
        RECT 50.165 50.025 52.775 50.055 ;
        RECT 50.165 47.970 50.790 50.025 ;
        RECT 50.165 47.940 52.525 47.970 ;
        RECT 45.255 47.770 52.525 47.940 ;
        RECT 45.255 47.740 47.865 47.770 ;
        RECT 50.165 47.740 52.525 47.770 ;
        RECT 45.255 47.535 45.425 47.740 ;
        RECT 45.225 47.475 45.455 47.535 ;
        RECT 45.130 46.475 45.550 47.475 ;
        RECT 45.225 45.035 45.455 46.475 ;
        RECT 45.255 44.830 45.425 45.035 ;
        RECT 46.180 44.830 47.220 47.740 ;
        RECT 47.915 47.475 48.145 47.535 ;
        RECT 49.885 47.475 50.115 47.535 ;
        RECT 47.850 46.475 48.210 47.475 ;
        RECT 49.820 46.475 50.180 47.475 ;
        RECT 47.915 45.035 48.145 46.475 ;
        RECT 49.885 45.035 50.115 46.475 ;
        RECT 50.765 44.830 51.805 47.740 ;
        RECT 52.575 46.095 52.805 47.535 ;
        RECT 52.480 45.095 52.900 46.095 ;
        RECT 52.575 45.035 52.805 45.095 ;
        RECT 45.255 44.600 47.865 44.830 ;
        RECT 50.165 44.600 52.525 44.830 ;
        RECT 53.225 44.345 53.930 53.970 ;
        RECT 59.190 52.020 59.885 55.000 ;
        RECT 60.415 54.530 60.875 54.760 ;
        RECT 61.205 54.530 61.665 54.760 ;
        RECT 61.995 54.530 62.455 54.760 ;
        RECT 62.785 54.530 63.245 54.760 ;
        RECT 60.135 53.885 60.365 54.325 ;
        RECT 60.070 53.385 60.430 53.885 ;
        RECT 60.135 53.325 60.365 53.385 ;
        RECT 60.575 53.120 60.755 54.530 ;
        RECT 61.325 54.525 61.505 54.530 ;
        RECT 60.925 53.325 61.155 54.325 ;
        RECT 61.330 53.125 61.495 54.525 ;
        RECT 61.715 54.265 61.945 54.325 ;
        RECT 61.650 53.765 62.010 54.265 ;
        RECT 61.715 53.325 61.945 53.765 ;
        RECT 61.325 53.120 61.505 53.125 ;
        RECT 62.150 53.120 62.330 54.530 ;
        RECT 62.505 53.325 62.735 54.325 ;
        RECT 62.910 53.120 63.090 54.530 ;
        RECT 63.295 53.885 63.525 54.325 ;
        RECT 63.230 53.385 63.590 53.885 ;
        RECT 63.295 53.325 63.525 53.385 ;
        RECT 60.415 52.890 60.875 53.120 ;
        RECT 61.205 52.890 61.665 53.120 ;
        RECT 61.995 52.890 62.455 53.120 ;
        RECT 62.785 52.890 63.245 53.120 ;
        RECT 59.210 51.960 59.865 52.020 ;
        RECT 60.415 51.745 60.665 52.890 ;
        RECT 60.415 51.475 61.065 51.745 ;
        RECT 60.415 50.565 60.665 51.475 ;
        RECT 57.545 50.315 60.665 50.565 ;
        RECT 56.175 49.490 56.580 49.550 ;
        RECT 56.155 46.465 56.600 49.490 ;
        RECT 57.545 48.640 57.795 50.315 ;
        RECT 61.205 50.075 61.455 52.890 ;
        RECT 61.995 51.130 62.245 52.890 ;
        RECT 61.600 50.860 62.245 51.130 ;
        RECT 60.325 49.825 61.455 50.075 ;
        RECT 61.995 50.075 62.245 50.860 ;
        RECT 62.785 50.565 63.035 52.890 ;
        RECT 63.815 52.090 64.555 55.000 ;
        RECT 68.725 54.235 102.145 55.160 ;
        RECT 63.835 52.030 64.535 52.090 ;
        RECT 62.785 50.315 65.925 50.565 ;
        RECT 61.995 49.825 63.145 50.075 ;
        RECT 57.335 48.410 57.795 48.640 ;
        RECT 57.055 48.190 57.285 48.250 ;
        RECT 56.990 47.790 57.350 48.190 ;
        RECT 57.055 47.250 57.285 47.790 ;
        RECT 57.845 47.710 58.075 48.250 ;
        RECT 57.780 47.310 58.140 47.710 ;
        RECT 57.845 47.250 58.075 47.310 ;
        RECT 57.335 46.860 57.795 47.090 ;
        RECT 58.585 46.465 59.270 49.550 ;
        RECT 60.325 48.640 60.575 49.825 ;
        RECT 60.115 48.410 60.575 48.640 ;
        RECT 59.835 47.710 60.065 48.250 ;
        RECT 60.625 48.190 60.855 48.250 ;
        RECT 60.560 47.790 60.920 48.190 ;
        RECT 59.770 47.310 60.130 47.710 ;
        RECT 59.835 47.250 60.065 47.310 ;
        RECT 60.625 47.250 60.855 47.790 ;
        RECT 60.115 46.860 60.575 47.090 ;
        RECT 60.125 46.780 60.565 46.860 ;
        RECT 61.370 46.465 62.055 49.565 ;
        RECT 62.895 48.640 63.145 49.825 ;
        RECT 62.895 48.410 63.355 48.640 ;
        RECT 62.615 48.190 62.845 48.250 ;
        RECT 62.550 47.790 62.910 48.190 ;
        RECT 62.615 47.250 62.845 47.790 ;
        RECT 63.405 47.710 63.635 48.250 ;
        RECT 63.340 47.310 63.700 47.710 ;
        RECT 63.405 47.250 63.635 47.310 ;
        RECT 62.895 46.860 63.355 47.090 ;
        RECT 64.190 46.465 64.875 49.525 ;
        RECT 65.675 48.640 65.925 50.315 ;
        RECT 66.890 49.500 67.270 49.560 ;
        RECT 65.675 48.410 66.135 48.640 ;
        RECT 65.395 47.710 65.625 48.250 ;
        RECT 66.185 48.190 66.415 48.250 ;
        RECT 66.120 47.790 66.480 48.190 ;
        RECT 65.330 47.310 65.690 47.710 ;
        RECT 65.395 47.250 65.625 47.310 ;
        RECT 66.185 47.250 66.415 47.790 ;
        RECT 65.675 46.860 66.135 47.090 ;
        RECT 65.685 46.780 66.125 46.860 ;
        RECT 66.870 46.465 67.290 49.500 ;
        RECT 56.145 45.835 67.290 46.465 ;
        RECT 29.190 43.775 30.355 43.805 ;
        RECT 44.010 43.705 53.930 44.345 ;
        RECT 44.030 43.655 53.930 43.705 ;
        RECT 44.030 43.645 44.780 43.655 ;
        RECT 53.225 43.640 53.930 43.655 ;
        RECT 53.245 43.580 53.910 43.640 ;
        RECT 42.585 43.250 42.975 43.310 ;
        RECT 42.565 43.230 42.995 43.250 ;
        RECT 26.530 43.210 42.995 43.230 ;
        RECT 26.445 43.160 42.995 43.210 ;
        RECT 26.445 43.150 54.010 43.160 ;
        RECT 26.425 42.790 54.010 43.150 ;
        RECT 26.425 42.770 42.995 42.790 ;
        RECT 26.425 40.075 26.925 42.770 ;
        RECT 27.575 42.355 33.535 42.385 ;
        RECT 35.855 42.355 41.815 42.385 ;
        RECT 27.325 42.185 41.815 42.355 ;
        RECT 27.325 42.155 33.535 42.185 ;
        RECT 35.855 42.155 41.815 42.185 ;
        RECT 27.325 41.995 27.495 42.155 ;
        RECT 27.295 41.935 27.525 41.995 ;
        RECT 33.585 41.935 33.815 41.995 ;
        RECT 35.575 41.935 35.805 41.995 ;
        RECT 27.200 41.615 27.620 41.935 ;
        RECT 27.295 40.995 27.525 41.615 ;
        RECT 33.520 41.435 33.880 41.935 ;
        RECT 35.510 41.435 35.870 41.935 ;
        RECT 33.585 40.995 33.815 41.435 ;
        RECT 35.575 40.995 35.805 41.435 ;
        RECT 41.865 41.375 42.095 41.995 ;
        RECT 41.770 41.055 42.190 41.375 ;
        RECT 41.865 40.995 42.095 41.055 ;
        RECT 27.320 40.835 27.495 40.995 ;
        RECT 27.320 40.805 33.535 40.835 ;
        RECT 35.855 40.805 41.815 40.835 ;
        RECT 27.320 40.635 41.815 40.805 ;
        RECT 27.320 40.605 33.535 40.635 ;
        RECT 35.855 40.605 41.815 40.635 ;
        RECT 42.565 40.075 42.995 42.770 ;
        RECT 26.425 40.005 42.995 40.075 ;
        RECT 44.070 40.005 44.855 42.790 ;
        RECT 45.505 42.155 47.665 42.385 ;
        RECT 45.225 41.935 45.455 41.995 ;
        RECT 45.130 41.435 45.550 41.935 ;
        RECT 47.715 41.555 47.945 41.995 ;
        RECT 45.225 40.995 45.455 41.435 ;
        RECT 47.650 41.055 48.010 41.555 ;
        RECT 47.715 40.995 47.945 41.055 ;
        RECT 45.515 40.835 46.415 40.855 ;
        RECT 45.505 40.605 47.665 40.835 ;
        RECT 45.515 40.535 46.415 40.605 ;
        RECT 48.470 40.005 49.535 42.790 ;
        RECT 50.365 42.160 52.525 42.390 ;
        RECT 50.085 41.940 50.315 42.000 ;
        RECT 52.575 41.940 52.805 42.000 ;
        RECT 50.020 41.440 50.380 41.940 ;
        RECT 52.480 41.440 52.900 41.940 ;
        RECT 50.085 41.000 50.315 41.440 ;
        RECT 52.575 41.000 52.805 41.440 ;
        RECT 50.375 40.840 51.275 40.865 ;
        RECT 50.365 40.610 52.525 40.840 ;
        RECT 50.375 40.545 51.275 40.610 ;
        RECT 53.275 40.005 54.000 42.790 ;
        RECT 26.425 39.635 54.070 40.005 ;
        RECT 26.425 39.315 42.995 39.635 ;
        RECT 26.425 36.505 26.925 39.315 ;
        RECT 27.325 38.775 33.535 38.805 ;
        RECT 35.855 38.775 41.815 38.805 ;
        RECT 27.325 38.605 41.815 38.775 ;
        RECT 27.325 38.575 33.535 38.605 ;
        RECT 35.855 38.575 41.815 38.605 ;
        RECT 27.325 38.415 27.495 38.575 ;
        RECT 27.295 38.355 27.525 38.415 ;
        RECT 27.200 38.035 27.620 38.355 ;
        RECT 27.295 37.415 27.525 38.035 ;
        RECT 33.585 37.975 33.815 38.415 ;
        RECT 35.575 37.975 35.805 38.415 ;
        RECT 33.520 37.475 33.880 37.975 ;
        RECT 35.510 37.475 35.870 37.975 ;
        RECT 41.865 37.740 42.095 38.415 ;
        RECT 33.585 37.415 33.815 37.475 ;
        RECT 35.575 37.415 35.805 37.475 ;
        RECT 41.770 37.420 42.190 37.740 ;
        RECT 41.865 37.415 42.095 37.420 ;
        RECT 27.325 37.255 27.495 37.415 ;
        RECT 27.325 37.225 33.535 37.255 ;
        RECT 35.855 37.225 41.815 37.255 ;
        RECT 27.325 37.055 41.815 37.225 ;
        RECT 27.325 37.025 33.535 37.055 ;
        RECT 35.855 37.025 41.815 37.055 ;
        RECT 42.565 36.505 42.995 39.315 ;
        RECT 26.425 35.745 42.995 36.505 ;
        RECT 26.425 32.850 26.925 35.745 ;
        RECT 27.575 35.195 33.535 35.225 ;
        RECT 35.855 35.195 42.065 35.225 ;
        RECT 27.575 35.025 42.065 35.195 ;
        RECT 27.575 34.995 33.535 35.025 ;
        RECT 35.855 34.995 42.065 35.025 ;
        RECT 41.895 34.835 42.065 34.995 ;
        RECT 27.295 34.775 27.525 34.835 ;
        RECT 27.200 34.455 27.620 34.775 ;
        RECT 27.295 33.835 27.525 34.455 ;
        RECT 33.585 34.395 33.815 34.835 ;
        RECT 35.575 34.395 35.805 34.835 ;
        RECT 41.865 34.775 42.095 34.835 ;
        RECT 41.770 34.455 42.190 34.775 ;
        RECT 33.520 33.895 33.880 34.395 ;
        RECT 35.510 33.895 35.870 34.395 ;
        RECT 33.585 33.835 33.815 33.895 ;
        RECT 35.575 33.835 35.805 33.895 ;
        RECT 41.865 33.835 42.095 34.455 ;
        RECT 41.895 33.675 42.065 33.835 ;
        RECT 27.575 33.645 33.535 33.675 ;
        RECT 35.855 33.645 42.065 33.675 ;
        RECT 27.575 33.475 42.065 33.645 ;
        RECT 27.575 33.445 33.535 33.475 ;
        RECT 35.855 33.445 42.065 33.475 ;
        RECT 42.565 32.850 42.995 35.745 ;
        RECT 26.425 32.090 42.995 32.850 ;
        RECT 26.425 29.365 26.925 32.090 ;
        RECT 27.575 31.615 33.535 31.645 ;
        RECT 35.855 31.615 42.065 31.645 ;
        RECT 27.575 31.445 42.065 31.615 ;
        RECT 27.575 31.415 33.535 31.445 ;
        RECT 35.855 31.415 42.065 31.445 ;
        RECT 41.895 31.255 42.065 31.415 ;
        RECT 27.295 30.635 27.525 31.255 ;
        RECT 33.585 30.815 33.815 31.255 ;
        RECT 35.575 30.815 35.805 31.255 ;
        RECT 41.865 31.195 42.095 31.255 ;
        RECT 41.770 30.875 42.190 31.195 ;
        RECT 27.200 30.315 27.620 30.635 ;
        RECT 33.520 30.315 33.880 30.815 ;
        RECT 35.510 30.315 35.870 30.815 ;
        RECT 27.295 30.255 27.525 30.315 ;
        RECT 33.585 30.255 33.815 30.315 ;
        RECT 35.575 30.255 35.805 30.315 ;
        RECT 41.865 30.255 42.095 30.875 ;
        RECT 41.895 30.095 42.065 30.255 ;
        RECT 27.575 30.065 33.535 30.095 ;
        RECT 35.855 30.065 42.065 30.095 ;
        RECT 27.575 29.895 42.065 30.065 ;
        RECT 27.575 29.865 33.535 29.895 ;
        RECT 35.855 29.865 42.065 29.895 ;
        RECT 42.565 29.365 42.995 32.090 ;
        RECT 26.425 28.650 42.995 29.365 ;
        RECT 26.445 28.605 42.995 28.650 ;
        RECT 26.445 28.590 26.905 28.605 ;
        RECT 42.565 28.600 42.995 28.605 ;
        RECT 42.585 28.540 42.975 28.600 ;
        RECT 68.725 11.985 69.395 54.235 ;
        RECT 70.765 53.455 72.045 53.485 ;
        RECT 73.725 53.455 75.155 53.485 ;
        RECT 76.670 53.455 78.100 53.485 ;
        RECT 79.585 53.455 81.015 53.485 ;
        RECT 70.535 51.350 72.265 53.455 ;
        RECT 73.495 51.350 75.225 53.455 ;
        RECT 76.455 51.350 78.185 53.455 ;
        RECT 79.415 51.350 81.145 53.455 ;
        RECT 70.765 51.325 72.045 51.350 ;
        RECT 73.725 51.325 75.155 51.350 ;
        RECT 76.670 51.325 78.100 51.350 ;
        RECT 79.585 51.325 81.015 51.350 ;
        RECT 82.830 49.675 102.115 54.235 ;
        RECT 83.015 48.600 100.625 48.830 ;
        RECT 83.015 40.500 83.245 48.600 ;
        RECT 83.805 48.380 84.035 48.440 ;
        RECT 83.740 46.380 84.100 48.380 ;
        RECT 82.950 38.500 83.310 40.500 ;
        RECT 83.015 38.280 83.245 38.500 ;
        RECT 83.805 38.440 84.035 46.380 ;
        RECT 84.595 40.500 84.825 48.600 ;
        RECT 85.385 48.380 85.615 48.440 ;
        RECT 85.320 46.380 85.680 48.380 ;
        RECT 84.530 38.500 84.890 40.500 ;
        RECT 84.595 38.280 84.825 38.500 ;
        RECT 85.385 38.440 85.615 46.380 ;
        RECT 86.175 40.500 86.405 48.600 ;
        RECT 86.965 48.380 87.195 48.440 ;
        RECT 86.900 46.380 87.260 48.380 ;
        RECT 86.110 38.500 86.470 40.500 ;
        RECT 86.175 38.280 86.405 38.500 ;
        RECT 86.965 38.440 87.195 46.380 ;
        RECT 87.755 40.500 87.985 48.600 ;
        RECT 88.545 48.380 88.775 48.440 ;
        RECT 88.480 46.380 88.840 48.380 ;
        RECT 87.690 38.500 88.050 40.500 ;
        RECT 87.755 38.280 87.985 38.500 ;
        RECT 88.545 38.440 88.775 46.380 ;
        RECT 89.335 40.500 89.565 48.600 ;
        RECT 90.125 48.385 90.355 48.440 ;
        RECT 90.060 46.385 90.420 48.385 ;
        RECT 89.270 38.500 89.630 40.500 ;
        RECT 89.335 38.280 89.565 38.500 ;
        RECT 90.125 38.440 90.355 46.385 ;
        RECT 90.915 40.500 91.145 48.600 ;
        RECT 91.705 48.380 91.935 48.440 ;
        RECT 91.640 46.380 92.000 48.380 ;
        RECT 90.850 38.500 91.210 40.500 ;
        RECT 90.915 38.280 91.145 38.500 ;
        RECT 91.705 38.440 91.935 46.380 ;
        RECT 92.495 40.500 92.725 48.600 ;
        RECT 93.285 48.380 93.515 48.440 ;
        RECT 93.220 46.380 93.580 48.380 ;
        RECT 92.430 38.500 92.790 40.500 ;
        RECT 92.495 38.280 92.725 38.500 ;
        RECT 93.285 38.440 93.515 46.380 ;
        RECT 94.075 40.500 94.305 48.600 ;
        RECT 94.865 48.380 95.095 48.440 ;
        RECT 94.800 46.380 95.160 48.380 ;
        RECT 94.010 38.500 94.370 40.500 ;
        RECT 94.075 38.280 94.305 38.500 ;
        RECT 94.865 38.440 95.095 46.380 ;
        RECT 95.655 40.500 95.885 48.600 ;
        RECT 96.445 48.380 96.675 48.440 ;
        RECT 96.380 46.380 96.740 48.380 ;
        RECT 95.590 38.500 95.950 40.500 ;
        RECT 95.655 38.280 95.885 38.500 ;
        RECT 96.445 38.440 96.675 46.380 ;
        RECT 97.235 40.500 97.465 48.600 ;
        RECT 98.025 48.380 98.255 48.440 ;
        RECT 97.960 46.380 98.320 48.380 ;
        RECT 97.170 38.500 97.530 40.500 ;
        RECT 97.235 38.280 97.465 38.500 ;
        RECT 98.025 38.440 98.255 46.380 ;
        RECT 98.815 40.500 99.045 48.600 ;
        RECT 99.605 48.380 99.835 48.440 ;
        RECT 99.540 46.380 99.900 48.380 ;
        RECT 98.750 38.500 99.110 40.500 ;
        RECT 98.815 38.280 99.045 38.500 ;
        RECT 99.605 38.440 99.835 46.380 ;
        RECT 100.395 40.500 100.625 48.600 ;
        RECT 101.340 48.685 102.115 49.675 ;
        RECT 101.340 47.440 102.030 48.685 ;
        RECT 100.330 38.500 100.690 40.500 ;
        RECT 100.395 38.280 100.625 38.500 ;
        RECT 83.015 38.050 100.625 38.280 ;
        RECT 101.255 37.425 102.030 47.440 ;
        RECT 121.785 40.870 123.125 40.900 ;
        RECT 106.565 40.820 120.185 40.835 ;
        RECT 106.550 40.785 120.510 40.820 ;
        RECT 105.945 40.725 120.510 40.785 ;
        RECT 100.770 37.395 102.030 37.425 ;
        RECT 82.295 36.420 102.030 37.395 ;
        RECT 91.665 36.215 102.030 36.420 ;
        RECT 72.185 35.960 73.615 35.985 ;
        RECT 75.150 35.960 76.580 35.985 ;
        RECT 78.070 35.960 79.500 35.985 ;
        RECT 70.535 33.990 70.785 35.960 ;
        RECT 70.485 32.495 70.835 33.990 ;
        RECT 72.015 33.855 73.745 35.960 ;
        RECT 74.975 33.855 76.705 35.960 ;
        RECT 77.935 33.855 79.665 35.960 ;
        RECT 80.895 35.915 81.145 35.960 ;
        RECT 83.415 35.915 84.395 35.930 ;
        RECT 86.345 35.915 87.325 35.930 ;
        RECT 89.275 35.915 90.255 35.930 ;
        RECT 80.840 33.915 81.200 35.915 ;
        RECT 83.405 35.685 84.405 35.915 ;
        RECT 86.335 35.685 87.335 35.915 ;
        RECT 89.265 35.685 90.265 35.915 ;
        RECT 83.415 35.670 84.395 35.685 ;
        RECT 86.345 35.670 87.325 35.685 ;
        RECT 89.275 35.670 90.255 35.685 ;
        RECT 83.015 35.210 83.245 35.635 ;
        RECT 84.565 35.210 86.175 35.635 ;
        RECT 87.495 35.620 87.770 35.635 ;
        RECT 88.830 35.620 89.105 35.635 ;
        RECT 87.495 35.605 87.775 35.620 ;
        RECT 88.820 35.605 89.105 35.620 ;
        RECT 87.495 35.210 89.105 35.605 ;
        RECT 90.425 35.210 90.655 35.635 ;
        RECT 80.895 33.855 81.145 33.915 ;
        RECT 72.185 33.825 73.615 33.855 ;
        RECT 75.150 33.825 76.580 33.855 ;
        RECT 78.070 33.825 79.500 33.855 ;
        RECT 72.160 32.665 73.540 32.695 ;
        RECT 75.170 32.665 76.550 32.695 ;
        RECT 78.115 32.665 79.495 32.695 ;
        RECT 70.535 30.560 70.785 32.495 ;
        RECT 72.015 30.560 73.745 32.665 ;
        RECT 74.975 30.560 76.705 32.665 ;
        RECT 77.935 30.560 79.665 32.665 ;
        RECT 72.160 30.535 73.540 30.560 ;
        RECT 75.170 30.535 76.550 30.560 ;
        RECT 78.115 30.535 79.495 30.560 ;
        RECT 80.795 30.535 81.245 32.695 ;
        RECT 80.895 30.530 81.145 30.535 ;
        RECT 83.015 28.285 90.655 35.210 ;
        RECT 92.535 31.860 97.690 32.835 ;
        RECT 93.735 31.165 95.285 31.170 ;
        RECT 96.715 31.165 98.265 31.195 ;
        RECT 93.620 29.060 95.400 31.165 ;
        RECT 96.530 29.060 98.415 31.165 ;
        RECT 93.735 29.035 95.285 29.060 ;
        RECT 83.015 26.160 90.720 28.285 ;
        RECT 83.015 26.110 86.175 26.160 ;
        RECT 83.015 25.675 83.245 26.110 ;
        RECT 84.565 25.675 86.175 26.110 ;
        RECT 87.495 25.745 89.105 26.160 ;
        RECT 87.495 25.690 87.775 25.745 ;
        RECT 88.820 25.690 89.105 25.745 ;
        RECT 90.360 25.735 90.720 26.160 ;
        RECT 87.495 25.675 87.770 25.690 ;
        RECT 88.830 25.675 89.105 25.690 ;
        RECT 90.425 25.675 90.655 25.735 ;
        RECT 83.415 25.625 84.395 25.640 ;
        RECT 86.345 25.625 87.325 25.640 ;
        RECT 89.275 25.625 90.255 25.640 ;
        RECT 83.405 25.395 84.405 25.625 ;
        RECT 86.335 25.395 87.335 25.625 ;
        RECT 89.265 25.395 90.265 25.625 ;
        RECT 83.415 25.380 84.395 25.395 ;
        RECT 86.345 25.380 87.325 25.395 ;
        RECT 89.275 25.380 90.255 25.395 ;
        RECT 83.415 23.605 84.395 23.620 ;
        RECT 86.345 23.605 87.325 23.620 ;
        RECT 89.275 23.605 90.255 23.620 ;
        RECT 83.405 23.375 84.405 23.605 ;
        RECT 86.335 23.375 87.335 23.605 ;
        RECT 89.265 23.375 90.265 23.605 ;
        RECT 83.415 23.360 84.395 23.375 ;
        RECT 86.345 23.360 87.325 23.375 ;
        RECT 89.275 23.360 90.255 23.375 ;
        RECT 70.705 15.170 72.085 15.195 ;
        RECT 73.700 15.170 75.080 15.195 ;
        RECT 76.615 15.170 77.995 15.195 ;
        RECT 79.620 15.170 81.000 15.195 ;
        RECT 70.535 13.065 72.265 15.170 ;
        RECT 73.495 13.065 75.225 15.170 ;
        RECT 76.455 13.065 78.185 15.170 ;
        RECT 79.415 13.065 81.145 15.170 ;
        RECT 83.015 13.365 83.245 23.325 ;
        RECT 84.565 13.365 86.175 23.325 ;
        RECT 87.495 13.365 89.105 23.325 ;
        RECT 90.425 15.925 90.655 23.325 ;
        RECT 90.360 13.425 90.720 15.925 ;
        RECT 90.425 13.365 90.655 13.425 ;
        RECT 83.415 13.315 84.395 13.330 ;
        RECT 86.345 13.315 87.325 13.330 ;
        RECT 89.275 13.315 90.255 13.330 ;
        RECT 83.405 13.085 84.405 13.315 ;
        RECT 86.335 13.085 87.335 13.315 ;
        RECT 89.265 13.085 90.265 13.315 ;
        RECT 83.415 13.070 84.395 13.085 ;
        RECT 86.345 13.070 87.325 13.085 ;
        RECT 89.275 13.070 90.255 13.085 ;
        RECT 70.705 13.035 72.085 13.065 ;
        RECT 73.700 13.035 75.080 13.065 ;
        RECT 76.615 13.035 77.995 13.065 ;
        RECT 79.620 13.035 81.000 13.065 ;
        RECT 93.520 13.035 93.970 15.195 ;
        RECT 95.050 13.065 96.880 15.170 ;
        RECT 95.265 13.035 96.815 13.065 ;
        RECT 97.960 13.035 98.415 15.195 ;
        RECT 100.445 11.985 102.030 36.215 ;
        RECT 105.925 40.110 120.510 40.725 ;
        RECT 121.785 40.490 134.235 40.870 ;
        RECT 121.785 40.170 134.225 40.490 ;
        RECT 105.925 29.850 107.570 40.110 ;
        RECT 114.975 39.755 118.675 39.770 ;
        RECT 108.685 39.525 118.685 39.755 ;
        RECT 114.975 39.510 118.675 39.525 ;
        RECT 108.295 39.045 108.525 39.475 ;
        RECT 108.295 37.060 108.600 39.045 ;
        RECT 118.845 37.060 119.075 39.475 ;
        RECT 119.525 39.045 120.480 40.110 ;
        RECT 121.785 39.115 123.125 40.170 ;
        RECT 123.720 39.755 127.115 39.770 ;
        RECT 123.720 39.525 128.590 39.755 ;
        RECT 123.720 39.510 127.115 39.525 ;
        RECT 123.720 39.275 123.950 39.510 ;
        RECT 128.360 39.275 128.590 39.525 ;
        RECT 108.295 35.635 119.075 37.060 ;
        RECT 108.220 33.735 119.075 35.635 ;
        RECT 108.220 30.635 108.600 33.735 ;
        RECT 118.845 33.560 119.075 33.735 ;
        RECT 118.845 30.945 119.170 33.560 ;
        RECT 108.295 30.515 108.525 30.635 ;
        RECT 108.695 30.465 112.395 30.480 ;
        RECT 108.685 30.235 118.685 30.465 ;
        RECT 108.695 30.220 112.395 30.235 ;
        RECT 105.925 28.945 118.675 29.850 ;
        RECT 118.835 29.185 119.170 30.945 ;
        RECT 105.925 17.985 107.570 28.945 ;
        RECT 108.295 28.935 108.525 28.945 ;
        RECT 108.695 28.505 112.395 28.520 ;
        RECT 108.685 28.275 118.685 28.505 ;
        RECT 108.695 28.260 112.395 28.275 ;
        RECT 108.295 28.040 108.525 28.250 ;
        RECT 108.220 27.725 108.600 28.040 ;
        RECT 108.220 26.425 108.595 27.725 ;
        RECT 108.295 25.995 108.595 26.425 ;
        RECT 118.830 27.180 119.170 29.185 ;
        RECT 118.830 25.995 119.165 27.180 ;
        RECT 108.295 25.955 119.165 25.995 ;
        RECT 108.295 24.325 119.075 25.955 ;
        RECT 108.215 22.670 119.075 24.325 ;
        RECT 108.215 19.325 108.595 22.670 ;
        RECT 118.830 19.715 119.075 22.670 ;
        RECT 119.495 21.585 120.510 39.045 ;
        RECT 121.790 38.860 123.120 39.115 ;
        RECT 121.770 25.155 123.140 38.860 ;
        RECT 123.720 38.650 128.590 39.275 ;
        RECT 123.720 26.855 123.950 38.650 ;
        RECT 128.360 38.515 128.590 38.650 ;
        RECT 125.195 38.465 128.145 38.480 ;
        RECT 124.155 38.235 128.155 38.465 ;
        RECT 125.195 38.220 128.145 38.235 ;
        RECT 129.120 37.715 134.225 40.170 ;
        RECT 124.355 36.740 134.225 37.715 ;
        RECT 124.165 36.225 127.865 36.240 ;
        RECT 124.155 35.995 132.655 36.225 ;
        RECT 124.165 35.980 127.865 35.995 ;
        RECT 128.945 34.935 132.645 34.950 ;
        RECT 124.155 34.705 132.655 34.935 ;
        RECT 128.945 34.690 132.645 34.705 ;
        RECT 124.165 33.645 127.865 33.660 ;
        RECT 124.155 33.415 132.655 33.645 ;
        RECT 124.165 33.400 127.865 33.415 ;
        RECT 128.945 32.355 132.645 32.370 ;
        RECT 124.155 32.125 132.655 32.355 ;
        RECT 128.945 32.110 132.645 32.125 ;
        RECT 124.165 31.065 127.865 31.080 ;
        RECT 124.155 30.835 132.655 31.065 ;
        RECT 124.165 30.820 127.865 30.835 ;
        RECT 128.945 29.775 132.645 29.790 ;
        RECT 124.155 29.545 132.655 29.775 ;
        RECT 128.945 29.530 132.645 29.545 ;
        RECT 124.165 28.485 127.865 28.500 ;
        RECT 124.155 28.255 132.655 28.485 ;
        RECT 124.165 28.240 127.865 28.255 ;
        RECT 128.950 27.195 132.650 27.210 ;
        RECT 124.155 26.965 132.655 27.195 ;
        RECT 128.950 26.950 132.650 26.965 ;
        RECT 123.645 26.015 124.025 26.855 ;
        RECT 123.720 25.955 123.950 26.015 ;
        RECT 132.860 25.955 133.090 35.965 ;
        RECT 133.490 28.005 134.225 36.740 ;
        RECT 133.510 26.670 134.205 28.005 ;
        RECT 124.165 25.905 127.865 25.920 ;
        RECT 124.155 25.675 132.655 25.905 ;
        RECT 124.165 25.660 127.865 25.675 ;
        RECT 133.495 25.155 134.230 26.670 ;
        RECT 121.730 22.675 134.230 25.155 ;
        RECT 121.730 22.315 134.235 22.675 ;
        RECT 134.120 21.585 134.555 21.615 ;
        RECT 119.495 20.265 134.585 21.585 ;
        RECT 119.525 20.235 134.585 20.265 ;
        RECT 120.040 20.220 134.585 20.235 ;
        RECT 118.845 19.650 119.075 19.715 ;
        RECT 108.295 19.265 108.525 19.325 ;
        RECT 118.845 19.295 119.080 19.650 ;
        RECT 118.845 19.265 119.075 19.295 ;
        RECT 114.975 19.215 118.675 19.230 ;
        RECT 123.340 19.215 127.040 19.230 ;
        RECT 108.685 18.985 118.685 19.215 ;
        RECT 123.330 18.985 133.330 19.215 ;
        RECT 114.975 18.970 118.675 18.985 ;
        RECT 123.340 18.970 127.040 18.985 ;
        RECT 119.525 17.985 120.480 18.780 ;
        RECT 122.940 18.575 123.170 18.935 ;
        RECT 105.925 16.370 121.565 17.985 ;
        RECT 122.840 16.370 123.170 18.575 ;
        RECT 133.490 16.370 133.720 18.935 ;
        RECT 105.925 16.230 121.625 16.370 ;
        RECT 105.925 16.165 121.565 16.230 ;
        RECT 105.935 15.975 121.565 16.165 ;
        RECT 105.935 15.500 121.525 15.975 ;
        RECT 105.965 12.015 106.670 15.500 ;
        RECT 107.480 14.795 120.050 15.025 ;
        RECT 107.200 14.575 107.430 14.635 ;
        RECT 107.135 13.575 107.495 14.575 ;
        RECT 68.725 11.315 102.030 11.985 ;
        RECT 68.735 11.265 102.030 11.315 ;
        RECT 68.735 11.235 69.395 11.265 ;
        RECT 93.120 11.245 93.370 11.265 ;
        RECT 100.770 11.210 102.030 11.265 ;
        RECT 105.065 10.175 106.690 12.015 ;
        RECT 105.965 8.950 106.670 10.175 ;
        RECT 107.200 9.635 107.430 13.575 ;
        RECT 107.665 9.490 108.250 14.795 ;
        RECT 108.490 10.695 108.720 14.635 ;
        RECT 108.425 9.695 108.785 10.695 ;
        RECT 108.490 9.635 108.720 9.695 ;
        RECT 107.490 9.475 108.250 9.490 ;
        RECT 108.990 9.475 109.575 14.795 ;
        RECT 109.780 14.575 110.010 14.635 ;
        RECT 109.715 13.575 110.075 14.575 ;
        RECT 109.780 9.635 110.010 13.575 ;
        RECT 110.270 9.475 110.855 14.795 ;
        RECT 111.070 10.695 111.300 14.635 ;
        RECT 111.005 9.695 111.365 10.695 ;
        RECT 111.070 9.635 111.300 9.695 ;
        RECT 111.570 9.475 112.155 14.795 ;
        RECT 112.360 14.575 112.590 14.635 ;
        RECT 112.295 13.575 112.655 14.575 ;
        RECT 112.360 9.635 112.590 13.575 ;
        RECT 112.810 9.475 113.395 14.795 ;
        RECT 113.650 10.695 113.880 14.635 ;
        RECT 113.585 9.695 113.945 10.695 ;
        RECT 113.650 9.635 113.880 9.695 ;
        RECT 114.135 9.475 114.720 14.795 ;
        RECT 114.940 14.575 115.170 14.635 ;
        RECT 114.875 13.575 115.235 14.575 ;
        RECT 114.940 9.635 115.170 13.575 ;
        RECT 115.405 9.475 115.990 14.795 ;
        RECT 116.230 10.695 116.460 14.635 ;
        RECT 116.165 9.695 116.525 10.695 ;
        RECT 116.230 9.635 116.460 9.695 ;
        RECT 116.715 9.475 117.300 14.795 ;
        RECT 117.520 14.575 117.750 14.635 ;
        RECT 117.455 13.575 117.815 14.575 ;
        RECT 117.520 9.635 117.750 13.575 ;
        RECT 118.015 9.475 118.600 14.795 ;
        RECT 118.810 10.695 119.040 14.635 ;
        RECT 118.745 9.695 119.105 10.695 ;
        RECT 118.810 9.635 119.040 9.695 ;
        RECT 119.300 9.475 119.885 14.795 ;
        RECT 120.100 14.575 120.330 14.635 ;
        RECT 120.035 13.575 120.395 14.575 ;
        RECT 120.100 9.635 120.330 13.575 ;
        RECT 107.480 9.245 120.050 9.475 ;
        RECT 120.885 9.300 121.525 15.500 ;
        RECT 122.840 14.075 133.720 16.370 ;
        RECT 122.940 13.045 133.720 14.075 ;
        RECT 122.940 9.975 123.170 13.045 ;
        RECT 133.490 9.975 133.720 13.045 ;
        RECT 123.340 9.925 127.040 9.935 ;
        RECT 123.330 9.695 133.330 9.925 ;
        RECT 123.340 9.675 127.040 9.695 ;
        RECT 134.100 9.300 134.575 20.220 ;
        RECT 107.490 9.230 108.250 9.245 ;
        RECT 120.885 8.950 134.575 9.300 ;
        RECT 105.965 8.315 134.575 8.950 ;
        RECT 105.965 8.285 134.555 8.315 ;
        RECT 105.965 8.250 121.535 8.285 ;
        RECT 105.965 8.220 106.670 8.250 ;
      LAYER met2 ;
        RECT 12.165 211.685 29.145 212.940 ;
        RECT 12.165 152.335 13.440 211.685 ;
        RECT 28.015 154.950 29.075 211.685 ;
        RECT 30.160 155.540 54.415 156.565 ;
        RECT 10.230 151.300 13.440 152.335 ;
        RECT 13.920 151.780 14.280 153.880 ;
        RECT 31.120 153.865 31.380 154.200 ;
        RECT 53.010 153.980 53.330 154.580 ;
        RECT 27.295 153.565 31.380 153.865 ;
        RECT 27.295 151.780 27.555 153.565 ;
        RECT 31.475 153.060 32.740 153.445 ;
        RECT 51.145 153.015 52.945 153.480 ;
        RECT 53.795 152.730 54.370 155.540 ;
        RECT 30.155 152.040 54.410 152.730 ;
        RECT 30.155 151.705 54.445 152.040 ;
        RECT 10.230 150.265 29.075 151.300 ;
        RECT 52.445 150.855 54.445 151.705 ;
        RECT 125.440 150.855 127.195 150.905 ;
        RECT 10.230 150.235 12.230 150.265 ;
        RECT 52.445 149.295 127.195 150.855 ;
        RECT 125.440 149.245 127.195 149.295 ;
        RECT 55.340 146.470 56.130 149.015 ;
        RECT 23.980 145.680 56.130 146.470 ;
        RECT 23.980 74.735 24.770 145.680 ;
        RECT 31.180 137.860 35.475 139.965 ;
        RECT 69.930 139.090 70.330 139.140 ;
        RECT 64.305 138.730 70.330 139.090 ;
        RECT 69.930 136.670 70.330 138.730 ;
        RECT 76.890 129.870 79.535 130.400 ;
        RECT 64.790 125.410 66.290 125.770 ;
        RECT 28.710 123.120 29.905 123.155 ;
        RECT 28.710 123.045 56.160 123.120 ;
        RECT 28.710 120.970 64.220 123.045 ;
        RECT 28.710 120.940 56.160 120.970 ;
        RECT 28.710 98.835 29.905 120.940 ;
        RECT 30.900 120.560 31.200 120.600 ;
        RECT 30.900 120.340 33.550 120.560 ;
        RECT 30.900 120.200 31.200 120.340 ;
        RECT 33.250 120.200 33.550 120.340 ;
        RECT 35.760 120.340 40.840 120.650 ;
        RECT 35.760 120.290 36.060 120.340 ;
        RECT 38.190 120.290 38.490 120.340 ;
        RECT 40.540 120.290 40.840 120.340 ;
        RECT 43.050 120.340 45.700 120.650 ;
        RECT 43.050 120.290 43.350 120.340 ;
        RECT 45.400 120.290 45.700 120.340 ;
        RECT 47.910 120.340 50.560 120.650 ;
        RECT 47.910 120.290 48.210 120.340 ;
        RECT 50.260 120.290 50.560 120.340 ;
        RECT 52.770 120.290 53.070 120.940 ;
        RECT 31.400 119.805 31.660 119.855 ;
        RECT 32.790 119.805 33.050 119.855 ;
        RECT 31.400 119.300 33.050 119.805 ;
        RECT 31.400 114.755 31.660 119.300 ;
        RECT 32.790 114.755 33.050 119.300 ;
        RECT 33.840 119.815 34.100 119.855 ;
        RECT 35.230 119.815 35.490 119.865 ;
        RECT 33.840 119.310 35.490 119.815 ;
        RECT 33.840 114.755 34.100 119.310 ;
        RECT 35.230 114.765 35.490 119.310 ;
        RECT 38.685 119.830 38.945 119.880 ;
        RECT 40.080 119.830 40.340 119.880 ;
        RECT 38.685 119.325 40.340 119.830 ;
        RECT 38.685 114.780 38.945 119.325 ;
        RECT 40.080 114.780 40.340 119.325 ;
        RECT 41.125 119.820 41.385 119.870 ;
        RECT 42.500 119.820 42.760 119.870 ;
        RECT 41.125 119.315 42.760 119.820 ;
        RECT 41.125 114.770 41.385 119.315 ;
        RECT 42.500 114.770 42.760 119.315 ;
        RECT 43.560 119.815 43.820 119.865 ;
        RECT 44.935 119.815 45.195 119.865 ;
        RECT 43.560 119.310 45.195 119.815 ;
        RECT 43.560 114.765 43.820 119.310 ;
        RECT 44.935 114.765 45.195 119.310 ;
        RECT 45.985 119.820 46.245 119.865 ;
        RECT 47.365 119.820 47.625 119.865 ;
        RECT 45.985 119.315 47.625 119.820 ;
        RECT 48.420 119.815 48.680 119.865 ;
        RECT 49.795 119.815 50.055 119.865 ;
        RECT 45.985 114.765 46.245 119.315 ;
        RECT 47.365 114.765 47.625 119.315 ;
        RECT 48.410 119.310 50.055 119.815 ;
        RECT 48.420 114.765 48.680 119.310 ;
        RECT 49.795 114.765 50.055 119.310 ;
        RECT 50.845 119.860 51.105 119.865 ;
        RECT 52.230 119.860 52.490 119.865 ;
        RECT 50.845 119.355 52.490 119.860 ;
        RECT 50.845 114.765 51.105 119.355 ;
        RECT 52.230 114.765 52.490 119.355 ;
        RECT 65.790 118.085 66.290 125.410 ;
        RECT 77.820 120.285 100.585 120.295 ;
        RECT 77.820 118.895 100.745 120.285 ;
        RECT 98.485 118.890 100.745 118.895 ;
        RECT 54.115 117.585 79.200 118.085 ;
        RECT 54.115 105.245 54.515 117.585 ;
        RECT 78.940 116.985 79.200 117.585 ;
        RECT 99.230 117.485 99.490 118.085 ;
        RECT 99.230 116.985 102.165 117.485 ;
        RECT 56.660 113.605 56.920 114.205 ;
        RECT 55.275 113.105 56.920 113.605 ;
        RECT 76.940 113.605 77.220 114.205 ;
        RECT 76.940 113.105 101.055 113.605 ;
        RECT 55.275 109.775 55.775 113.105 ;
        RECT 56.760 110.810 75.630 111.830 ;
        RECT 80.735 110.680 100.205 111.955 ;
        RECT 55.275 109.725 56.045 109.775 ;
        RECT 100.555 109.725 101.055 113.105 ;
        RECT 55.275 109.225 79.200 109.725 ;
        RECT 55.545 109.175 56.045 109.225 ;
        RECT 56.695 105.245 56.955 105.845 ;
        RECT 54.115 104.745 56.955 105.245 ;
        RECT 56.395 103.430 75.145 103.965 ;
        RECT 75.525 101.455 75.905 109.225 ;
        RECT 77.650 105.985 78.430 108.890 ;
        RECT 78.940 108.625 79.200 109.225 ;
        RECT 99.230 109.225 101.055 109.725 ;
        RECT 99.230 108.625 99.490 109.225 ;
        RECT 99.805 105.985 100.740 108.810 ;
        RECT 76.985 105.245 77.245 105.845 ;
        RECT 77.650 105.755 100.740 105.985 ;
        RECT 77.685 105.500 100.740 105.755 ;
        RECT 100.635 105.245 101.135 105.295 ;
        RECT 101.665 105.245 102.165 116.985 ;
        RECT 76.985 104.745 102.165 105.245 ;
        RECT 100.635 104.695 101.135 104.745 ;
        RECT 75.525 101.075 104.935 101.455 ;
        RECT 30.900 98.485 31.200 100.300 ;
        RECT 33.330 100.220 33.630 100.270 ;
        RECT 35.680 100.220 35.980 100.270 ;
        RECT 33.330 99.910 35.980 100.220 ;
        RECT 30.845 97.885 31.230 98.485 ;
        RECT 26.365 97.310 26.865 97.360 ;
        RECT 38.110 97.310 38.410 100.270 ;
        RECT 40.620 100.220 40.920 100.270 ;
        RECT 42.970 100.220 43.270 100.270 ;
        RECT 40.620 99.910 43.270 100.220 ;
        RECT 45.480 100.220 45.780 100.270 ;
        RECT 47.830 100.220 48.130 100.270 ;
        RECT 45.480 99.910 48.130 100.220 ;
        RECT 50.340 100.220 50.640 100.270 ;
        RECT 52.690 100.220 52.990 100.270 ;
        RECT 50.340 99.910 52.990 100.220 ;
        RECT 26.365 97.050 38.410 97.310 ;
        RECT 26.365 96.875 26.865 97.050 ;
        RECT 31.745 91.085 32.005 97.050 ;
        RECT 46.750 95.385 51.750 95.765 ;
        RECT 57.530 95.385 62.530 95.765 ;
        RECT 31.710 87.145 32.030 88.245 ;
        RECT 23.980 74.375 47.100 74.735 ;
        RECT 23.980 60.470 24.770 74.375 ;
        RECT 40.270 73.645 41.230 73.995 ;
        RECT 41.745 73.645 42.005 73.980 ;
        RECT 40.270 73.245 42.005 73.645 ;
        RECT 52.035 73.665 52.295 95.245 ;
        RECT 99.075 92.145 99.395 95.245 ;
        RECT 104.555 93.590 104.935 101.075 ;
        RECT 107.015 93.610 107.515 94.030 ;
        RECT 105.175 88.450 105.455 93.550 ;
        RECT 57.155 85.265 57.475 88.365 ;
        RECT 107.695 88.240 107.975 93.340 ;
        RECT 57.155 80.125 57.475 83.225 ;
        RECT 77.475 80.625 77.735 87.865 ;
        RECT 78.815 80.625 79.075 87.865 ;
        RECT 77.475 73.665 77.735 74.300 ;
        RECT 78.815 73.665 79.075 74.300 ;
        RECT 99.075 74.050 99.395 76.345 ;
        RECT 99.025 73.890 99.445 74.050 ;
        RECT 52.035 73.245 107.650 73.665 ;
        RECT 40.270 72.370 41.230 73.245 ;
        RECT 107.630 72.400 110.265 72.405 ;
        RECT 107.565 72.370 110.265 72.400 ;
        RECT 40.270 72.200 110.270 72.370 ;
        RECT 40.280 71.160 110.270 72.200 ;
        RECT 39.805 69.905 110.270 71.160 ;
        RECT 107.565 69.895 110.270 69.905 ;
        RECT 107.630 69.850 110.270 69.895 ;
        RECT 107.630 69.845 110.265 69.850 ;
        RECT 47.955 64.170 50.625 65.345 ;
        RECT 39.000 63.620 54.065 64.170 ;
        RECT 39.000 63.365 53.890 63.620 ;
        RECT 39.000 62.545 53.895 63.365 ;
        RECT 40.320 60.625 40.580 62.545 ;
        RECT 23.980 60.110 44.220 60.470 ;
        RECT 29.180 58.755 50.375 59.895 ;
        RECT 29.180 55.920 29.915 58.755 ;
        RECT 30.255 55.810 30.610 57.790 ;
        RECT 50.610 56.070 50.870 61.605 ;
        RECT 48.850 55.810 50.870 56.070 ;
        RECT 26.365 55.625 26.865 55.675 ;
        RECT 26.365 55.265 35.675 55.625 ;
        RECT 26.365 55.215 26.865 55.265 ;
        RECT 29.200 54.150 48.560 54.830 ;
        RECT 30.850 51.580 31.170 52.860 ;
        RECT 34.460 49.800 34.925 51.020 ;
        RECT 38.220 50.380 38.540 51.660 ;
        RECT 21.825 49.595 22.490 49.645 ;
        RECT 21.825 49.590 28.420 49.595 ;
        RECT 31.175 49.590 31.675 49.640 ;
        RECT 35.855 49.590 36.355 49.640 ;
        RECT 21.825 49.090 36.355 49.590 ;
        RECT 21.825 49.040 22.490 49.090 ;
        RECT 31.175 49.040 31.675 49.090 ;
        RECT 35.855 49.040 36.355 49.090 ;
        RECT 19.625 48.840 20.290 48.890 ;
        RECT 33.035 48.840 33.535 48.890 ;
        RECT 37.745 48.840 38.245 48.890 ;
        RECT 19.625 48.340 38.245 48.840 ;
        RECT 19.625 48.290 20.290 48.340 ;
        RECT 33.035 48.290 33.535 48.340 ;
        RECT 37.745 48.290 38.245 48.340 ;
        RECT 30.850 45.170 31.170 46.450 ;
        RECT 38.220 46.375 38.540 47.650 ;
        RECT 38.935 44.405 39.710 54.150 ;
        RECT 29.350 43.785 39.800 44.405 ;
        RECT 44.060 44.365 44.750 54.150 ;
        RECT 48.850 53.910 49.180 55.810 ;
        RECT 51.420 53.980 53.895 62.545 ;
        RECT 61.745 55.635 64.470 60.555 ;
        RECT 66.620 56.310 103.890 56.990 ;
        RECT 59.400 55.620 65.020 55.635 ;
        RECT 59.240 54.980 65.020 55.620 ;
        RECT 47.900 53.650 50.130 53.910 ;
        RECT 45.180 50.470 45.500 51.570 ;
        RECT 45.180 46.425 45.500 47.525 ;
        RECT 47.900 46.425 48.160 53.650 ;
        RECT 49.870 46.425 50.130 53.650 ;
        RECT 52.530 51.850 52.850 52.950 ;
        RECT 52.530 45.045 52.850 46.145 ;
        RECT 53.275 44.365 53.880 53.980 ;
        RECT 59.240 51.970 59.835 54.980 ;
        RECT 56.830 51.130 57.330 51.260 ;
        RECT 60.120 51.130 60.380 53.935 ;
        RECT 61.700 53.715 61.960 54.980 ;
        RECT 60.655 51.745 61.030 51.775 ;
        RECT 63.280 51.745 63.540 53.935 ;
        RECT 63.865 52.040 64.505 54.980 ;
        RECT 66.620 51.745 67.365 56.310 ;
        RECT 101.455 55.210 102.065 55.250 ;
        RECT 60.655 51.475 67.365 51.745 ;
        RECT 60.655 51.445 61.030 51.475 ;
        RECT 61.605 51.130 61.970 51.160 ;
        RECT 56.830 50.860 61.970 51.130 ;
        RECT 56.830 50.810 57.330 50.860 ;
        RECT 56.205 46.485 56.550 49.540 ;
        RECT 60.610 48.245 60.870 50.860 ;
        RECT 61.605 50.830 61.970 50.860 ;
        RECT 57.235 48.240 60.870 48.245 ;
        RECT 57.040 47.985 60.870 48.240 ;
        RECT 57.040 47.740 57.300 47.985 ;
        RECT 57.830 47.540 58.090 47.760 ;
        RECT 59.820 47.540 60.080 47.760 ;
        RECT 60.610 47.740 60.870 47.985 ;
        RECT 62.600 48.240 62.860 51.475 ;
        RECT 66.620 51.465 67.365 51.475 ;
        RECT 68.775 54.270 102.065 55.210 ;
        RECT 62.600 47.980 66.430 48.240 ;
        RECT 62.600 47.740 62.860 47.980 ;
        RECT 57.830 47.310 60.080 47.540 ;
        RECT 57.830 46.485 58.090 47.310 ;
        RECT 59.820 47.260 60.080 47.310 ;
        RECT 63.390 47.490 63.650 47.760 ;
        RECT 65.380 47.490 65.640 47.760 ;
        RECT 66.170 47.740 66.430 47.980 ;
        RECT 63.390 47.260 65.640 47.490 ;
        RECT 60.175 46.730 60.515 47.110 ;
        RECT 63.390 46.485 63.650 47.260 ;
        RECT 65.735 46.730 66.075 47.110 ;
        RECT 66.920 46.485 67.240 49.550 ;
        RECT 56.205 46.385 67.240 46.485 ;
        RECT 56.205 46.355 67.230 46.385 ;
        RECT 56.150 45.815 67.230 46.355 ;
        RECT 44.060 43.655 53.880 44.365 ;
        RECT 44.105 43.635 53.880 43.655 ;
        RECT 53.275 43.590 53.880 43.635 ;
        RECT 42.615 43.250 42.945 43.300 ;
        RECT 26.590 43.200 42.945 43.250 ;
        RECT 26.475 43.180 42.945 43.200 ;
        RECT 26.475 42.830 53.950 43.180 ;
        RECT 56.185 42.830 58.545 45.815 ;
        RECT 26.475 42.770 58.545 42.830 ;
        RECT 26.475 42.750 42.945 42.770 ;
        RECT 22.640 42.645 23.515 42.695 ;
        RECT 26.475 42.645 26.875 42.750 ;
        RECT 22.640 40.645 26.875 42.645 ;
        RECT 27.250 41.565 27.570 41.985 ;
        RECT 33.570 41.385 33.830 42.750 ;
        RECT 35.560 41.385 35.820 42.750 ;
        RECT 41.820 41.005 42.140 41.425 ;
        RECT 22.640 40.595 23.515 40.645 ;
        RECT 26.475 40.095 26.875 40.645 ;
        RECT 42.615 40.095 42.945 42.750 ;
        RECT 26.475 40.025 42.945 40.095 ;
        RECT 44.120 40.025 44.805 42.770 ;
        RECT 45.180 41.385 45.500 41.985 ;
        RECT 45.565 40.485 46.365 40.905 ;
        RECT 47.700 40.025 47.960 41.605 ;
        RECT 48.520 40.025 49.485 42.770 ;
        RECT 50.070 41.390 50.330 42.770 ;
        RECT 52.530 41.390 52.850 41.990 ;
        RECT 50.425 40.495 51.225 40.915 ;
        RECT 53.325 40.470 58.545 42.770 ;
        RECT 53.325 40.025 53.950 40.470 ;
        RECT 26.475 39.615 54.010 40.025 ;
        RECT 26.475 39.295 42.945 39.615 ;
        RECT 26.475 36.525 26.875 39.295 ;
        RECT 27.250 37.985 27.570 38.405 ;
        RECT 33.570 36.525 33.830 38.025 ;
        RECT 35.560 36.525 35.820 38.025 ;
        RECT 41.820 37.370 42.140 37.790 ;
        RECT 42.615 36.525 42.945 39.295 ;
        RECT 26.475 35.725 42.945 36.525 ;
        RECT 26.475 32.870 26.875 35.725 ;
        RECT 27.250 34.405 27.570 34.825 ;
        RECT 33.570 32.870 33.830 34.445 ;
        RECT 35.560 32.870 35.820 34.445 ;
        RECT 41.820 34.405 42.140 34.825 ;
        RECT 42.615 32.870 42.945 35.725 ;
        RECT 26.475 32.070 42.945 32.870 ;
        RECT 26.475 29.385 26.875 32.070 ;
        RECT 27.250 30.265 27.570 30.685 ;
        RECT 33.570 29.385 33.830 30.865 ;
        RECT 35.560 29.385 35.820 30.865 ;
        RECT 41.820 30.825 42.140 31.245 ;
        RECT 42.615 29.385 42.945 32.070 ;
        RECT 26.475 29.125 42.945 29.385 ;
        RECT 26.360 28.585 42.945 29.125 ;
        RECT 42.615 28.550 42.945 28.585 ;
        RECT 68.775 12.030 69.345 54.270 ;
        RECT 82.880 49.625 102.065 54.270 ;
        RECT 101.455 48.635 102.065 49.625 ;
        RECT 90.110 48.430 90.370 48.435 ;
        RECT 103.210 48.430 103.890 56.310 ;
        RECT 80.665 47.750 103.890 48.430 ;
        RECT 80.665 33.865 81.370 47.750 ;
        RECT 83.790 46.330 84.050 47.750 ;
        RECT 85.370 46.330 85.630 47.750 ;
        RECT 86.950 46.330 87.210 47.750 ;
        RECT 88.530 46.330 88.790 47.750 ;
        RECT 90.110 46.335 90.370 47.750 ;
        RECT 91.690 46.330 91.950 47.750 ;
        RECT 93.270 46.330 93.530 47.750 ;
        RECT 94.850 46.330 95.110 47.750 ;
        RECT 96.430 46.330 96.690 47.750 ;
        RECT 98.010 46.330 98.270 47.750 ;
        RECT 99.590 46.330 99.850 47.750 ;
        RECT 83.000 39.130 83.260 40.550 ;
        RECT 84.580 39.130 84.840 40.550 ;
        RECT 86.160 39.130 86.420 40.550 ;
        RECT 87.740 39.130 88.000 40.550 ;
        RECT 89.320 39.130 89.580 40.550 ;
        RECT 90.900 39.130 91.160 40.550 ;
        RECT 92.480 39.130 92.740 40.550 ;
        RECT 94.060 39.130 94.320 40.550 ;
        RECT 95.640 39.130 95.900 40.550 ;
        RECT 97.220 39.130 97.480 40.550 ;
        RECT 98.800 39.130 99.060 40.550 ;
        RECT 100.380 39.130 100.640 40.550 ;
        RECT 83.000 38.450 100.640 39.130 ;
        RECT 83.000 35.980 83.260 38.450 ;
        RECT 101.305 37.270 101.915 47.490 ;
        RECT 106.600 40.775 120.460 40.870 ;
        RECT 91.715 36.915 101.915 37.270 ;
        RECT 105.975 40.060 120.460 40.775 ;
        RECT 121.975 40.845 134.335 40.890 ;
        RECT 121.975 40.390 134.665 40.845 ;
        RECT 121.975 40.150 134.335 40.390 ;
        RECT 91.715 36.165 101.920 36.915 ;
        RECT 83.000 35.620 84.405 35.980 ;
        RECT 86.335 35.620 90.205 35.980 ;
        RECT 100.495 32.855 101.920 36.165 ;
        RECT 80.845 31.000 81.195 32.745 ;
        RECT 92.595 31.840 101.920 32.855 ;
        RECT 97.480 31.835 101.920 31.840 ;
        RECT 80.840 23.670 81.200 31.000 ;
        RECT 90.410 25.965 90.670 28.335 ;
        RECT 90.410 25.705 92.300 25.965 ;
        RECT 89.325 25.690 90.205 25.705 ;
        RECT 83.465 25.330 87.375 25.690 ;
        RECT 89.265 25.330 90.225 25.690 ;
        RECT 89.325 25.315 90.205 25.330 ;
        RECT 80.840 23.310 84.440 23.670 ;
        RECT 86.295 23.310 90.205 23.670 ;
        RECT 89.325 13.380 90.205 13.395 ;
        RECT 83.465 13.020 87.355 13.380 ;
        RECT 89.265 13.020 90.205 13.380 ;
        RECT 89.325 13.005 90.205 13.020 ;
        RECT 68.750 11.970 80.215 12.030 ;
        RECT 68.035 11.265 82.730 11.970 ;
        RECT 84.480 11.265 90.035 11.970 ;
        RECT 68.750 10.855 80.215 11.265 ;
        RECT 58.890 3.390 59.790 3.440 ;
        RECT 90.410 3.390 90.670 15.975 ;
        RECT 91.045 11.265 91.610 11.970 ;
        RECT 58.840 3.130 90.670 3.390 ;
        RECT 58.890 3.005 59.790 3.130 ;
        RECT 78.210 2.275 79.110 2.325 ;
        RECT 92.040 2.275 92.300 25.705 ;
        RECT 93.570 12.985 93.920 15.245 ;
        RECT 98.010 12.985 98.365 15.245 ;
        RECT 100.495 11.950 101.920 31.835 ;
        RECT 105.975 18.005 107.520 40.060 ;
        RECT 115.025 39.460 127.065 39.820 ;
        RECT 108.270 24.375 108.550 35.685 ;
        RECT 108.745 30.170 112.345 30.530 ;
        RECT 108.745 28.570 109.585 30.170 ;
        RECT 109.895 29.810 118.605 29.840 ;
        RECT 119.545 29.810 120.460 39.095 ;
        RECT 109.895 28.975 120.460 29.810 ;
        RECT 109.895 28.925 118.605 28.975 ;
        RECT 108.745 28.210 112.345 28.570 ;
        RECT 108.265 24.310 108.550 24.375 ;
        RECT 108.265 19.275 108.545 24.310 ;
        RECT 119.545 21.605 120.460 28.975 ;
        RECT 121.820 37.735 123.090 38.910 ;
        RECT 125.245 38.170 128.095 38.530 ;
        RECT 127.050 37.735 128.095 38.170 ;
        RECT 129.180 38.035 134.335 40.150 ;
        RECT 129.180 37.735 134.175 38.035 ;
        RECT 121.820 36.720 134.175 37.735 ;
        RECT 121.820 25.175 123.090 36.720 ;
        RECT 126.760 36.290 127.815 36.720 ;
        RECT 124.215 35.930 127.815 36.290 ;
        RECT 124.215 33.710 124.950 35.930 ;
        RECT 128.995 34.860 132.595 35.000 ;
        RECT 128.995 34.640 132.600 34.860 ;
        RECT 124.215 33.350 127.815 33.710 ;
        RECT 124.215 31.130 124.950 33.350 ;
        RECT 131.740 32.420 132.600 34.640 ;
        RECT 128.995 32.060 132.600 32.420 ;
        RECT 124.215 30.770 127.815 31.130 ;
        RECT 124.215 28.550 124.950 30.770 ;
        RECT 131.740 29.840 132.600 32.060 ;
        RECT 128.995 29.480 132.600 29.840 ;
        RECT 124.215 28.190 127.815 28.550 ;
        RECT 123.695 25.965 123.975 26.905 ;
        RECT 124.215 25.970 124.950 28.190 ;
        RECT 131.740 27.675 132.600 29.480 ;
        RECT 133.540 27.955 134.175 36.720 ;
        RECT 136.170 27.675 137.070 27.725 ;
        RECT 131.740 27.260 137.070 27.675 ;
        RECT 129.000 26.900 137.070 27.260 ;
        RECT 136.170 26.850 137.070 26.900 ;
        RECT 124.215 25.610 127.815 25.970 ;
        RECT 124.215 25.175 124.950 25.610 ;
        RECT 133.545 25.175 134.180 26.720 ;
        RECT 121.790 22.410 134.180 25.175 ;
        RECT 121.790 22.295 134.175 22.410 ;
        RECT 119.545 20.215 134.525 21.605 ;
        RECT 120.100 20.200 134.525 20.215 ;
        RECT 115.025 18.920 126.990 19.280 ;
        RECT 105.565 16.295 105.835 16.300 ;
        RECT 105.975 16.295 121.505 18.005 ;
        RECT 105.565 15.955 121.505 16.295 ;
        RECT 105.565 15.480 121.475 15.955 ;
        RECT 107.185 14.625 107.565 15.480 ;
        RECT 109.770 14.625 110.230 15.480 ;
        RECT 112.190 14.625 112.650 15.480 ;
        RECT 114.900 14.625 115.355 15.480 ;
        RECT 117.470 14.625 117.925 15.480 ;
        RECT 120.055 14.625 120.510 15.480 ;
        RECT 107.185 14.570 120.510 14.625 ;
        RECT 107.185 14.365 120.345 14.570 ;
        RECT 107.185 13.525 107.445 14.365 ;
        RECT 109.765 13.525 110.025 14.365 ;
        RECT 112.345 13.525 112.605 14.365 ;
        RECT 114.925 13.525 115.185 14.365 ;
        RECT 117.505 13.525 117.765 14.365 ;
        RECT 120.085 13.525 120.345 14.365 ;
        RECT 93.120 11.245 101.920 11.950 ;
        RECT 93.520 9.540 93.970 10.485 ;
        RECT 105.115 10.125 106.640 12.065 ;
        RECT 108.475 9.990 108.735 10.745 ;
        RECT 111.055 9.990 111.315 10.745 ;
        RECT 113.635 9.990 113.895 10.745 ;
        RECT 116.215 9.990 116.475 10.745 ;
        RECT 118.795 9.990 119.055 10.745 ;
        RECT 120.935 10.135 121.475 15.480 ;
        RECT 122.890 14.025 123.210 18.625 ;
        RECT 108.475 9.630 127.015 9.990 ;
        RECT 93.520 9.180 108.195 9.540 ;
        RECT 97.530 3.400 98.435 9.180 ;
        RECT 120.935 8.970 121.475 9.370 ;
        RECT 106.075 8.230 121.475 8.970 ;
        RECT 121.715 7.090 122.375 9.630 ;
        RECT 123.390 9.625 126.990 9.630 ;
        RECT 134.150 9.325 134.525 20.200 ;
        RECT 132.395 9.320 134.525 9.325 ;
        RECT 122.745 8.265 134.525 9.320 ;
        RECT 78.210 2.015 92.300 2.275 ;
        RECT 78.210 1.925 79.110 2.015 ;
      LAYER met3 ;
        RECT 57.220 186.135 89.080 213.910 ;
        RECT 91.700 186.135 123.560 213.920 ;
        RECT 57.220 183.520 123.560 186.135 ;
        RECT 57.220 183.510 93.400 183.520 ;
        RECT 86.725 181.630 93.400 183.510 ;
        RECT 57.215 181.620 93.400 181.630 ;
        RECT 57.215 179.550 123.555 181.620 ;
        RECT 52.960 154.005 53.465 154.560 ;
        RECT 10.180 150.260 12.280 152.310 ;
        RECT 13.870 151.805 14.330 153.855 ;
        RECT 57.215 153.455 89.075 179.550 ;
        RECT 31.425 153.085 32.790 153.420 ;
        RECT 13.920 149.655 14.280 151.805 ;
        RECT 28.420 151.165 29.100 151.190 ;
        RECT 31.425 151.165 31.820 153.085 ;
        RECT 51.095 153.040 89.075 153.455 ;
        RECT 57.215 151.230 89.075 153.040 ;
        RECT 91.695 151.220 123.555 179.550 ;
        RECT 28.420 150.780 31.820 151.165 ;
        RECT 28.420 150.755 29.100 150.780 ;
        RECT 13.845 67.800 14.345 149.655 ;
        RECT 125.390 149.270 127.245 150.880 ;
        RECT 55.290 147.970 56.180 148.990 ;
        RECT 31.130 137.885 35.525 139.940 ;
        RECT 76.840 129.895 79.585 130.375 ;
        RECT 27.450 120.225 31.250 120.575 ;
        RECT 76.890 113.130 77.270 129.895 ;
        RECT 98.435 120.250 100.795 120.260 ;
        RECT 110.320 120.250 139.680 135.540 ;
        RECT 98.435 118.950 139.680 120.250 ;
        RECT 98.435 118.915 100.795 118.950 ;
        RECT 55.495 109.200 56.095 109.750 ;
        RECT 110.320 107.640 139.680 118.950 ;
        RECT 100.585 104.720 101.185 105.270 ;
        RECT 135.505 104.610 139.160 107.640 ;
        RECT 30.795 97.910 31.280 98.460 ;
        RECT 26.315 96.900 26.915 97.335 ;
        RECT 46.700 95.410 62.580 95.740 ;
        RECT 99.025 92.170 99.445 95.220 ;
        RECT 105.125 93.635 107.565 94.040 ;
        RECT 105.125 93.630 107.135 93.635 ;
        RECT 105.125 88.475 105.505 93.630 ;
        RECT 110.320 93.315 139.680 104.610 ;
        RECT 107.645 92.815 139.680 93.315 ;
        RECT 31.660 87.170 32.080 88.220 ;
        RECT 57.105 85.290 57.525 88.340 ;
        RECT 107.645 88.265 108.025 92.815 ;
        RECT 57.105 80.150 57.525 83.200 ;
        RECT 110.320 76.710 139.680 92.815 ;
        RECT 99.025 73.845 99.445 76.320 ;
        RECT 107.580 72.345 110.315 72.380 ;
        RECT 107.580 69.875 110.320 72.345 ;
        RECT 107.580 69.870 110.315 69.875 ;
        RECT 13.845 67.300 57.330 67.800 ;
        RECT 47.905 64.610 50.675 65.320 ;
        RECT 30.205 56.330 30.660 57.765 ;
        RECT 30.205 55.835 34.975 56.330 ;
        RECT 30.215 55.830 34.975 55.835 ;
        RECT 26.315 55.240 26.915 55.650 ;
        RECT 30.800 51.605 31.220 52.835 ;
        RECT 34.410 49.825 34.975 55.830 ;
        RECT 43.805 52.605 52.900 52.925 ;
        RECT 38.170 50.905 38.590 51.635 ;
        RECT 38.170 50.405 39.905 50.905 ;
        RECT 21.775 49.065 22.540 49.620 ;
        RECT 19.575 48.315 20.340 48.865 ;
        RECT 30.800 45.695 31.220 46.425 ;
        RECT 38.170 46.400 38.590 47.625 ;
        RECT 39.405 45.695 39.905 50.405 ;
        RECT 43.805 47.500 44.125 52.605 ;
        RECT 52.480 51.875 52.900 52.605 ;
        RECT 45.130 50.495 45.550 51.545 ;
        RECT 56.830 51.235 57.330 67.300 ;
        RECT 61.695 59.605 64.520 60.530 ;
        RECT 56.780 50.835 57.380 51.235 ;
        RECT 43.805 47.180 45.550 47.500 ;
        RECT 30.800 45.195 39.905 45.695 ;
        RECT 22.590 42.645 23.565 42.670 ;
        RECT 14.310 40.645 23.565 42.645 ;
        RECT 27.195 41.590 27.935 41.960 ;
        RECT 30.800 41.940 31.220 45.195 ;
        RECT 38.165 43.375 38.595 43.695 ;
        RECT 30.755 41.610 31.270 41.940 ;
        RECT 38.215 41.275 38.545 43.375 ;
        RECT 45.130 41.410 45.550 47.180 ;
        RECT 52.480 45.070 52.900 46.120 ;
        RECT 52.480 41.415 52.900 42.200 ;
        RECT 41.770 41.275 42.190 41.400 ;
        RECT 22.590 40.620 23.565 40.645 ;
        RECT 25.965 40.930 42.190 41.275 ;
        RECT 25.965 38.380 26.335 40.930 ;
        RECT 45.515 40.510 46.415 40.880 ;
        RECT 50.375 40.520 51.275 40.890 ;
        RECT 50.375 38.385 50.695 40.520 ;
        RECT 43.535 38.380 50.695 38.385 ;
        RECT 25.965 38.065 50.695 38.380 ;
        RECT 25.965 38.010 27.830 38.065 ;
        RECT 25.965 30.660 26.335 38.010 ;
        RECT 41.440 37.395 42.190 37.765 ;
        RECT 43.550 34.800 43.920 38.065 ;
        RECT 27.200 34.430 27.900 34.800 ;
        RECT 41.770 34.430 43.920 34.800 ;
        RECT 41.530 30.850 42.215 31.220 ;
        RECT 25.965 30.290 27.620 30.660 ;
        RECT 27.410 12.010 29.235 12.035 ;
        RECT 14.925 10.175 29.240 12.010 ;
        RECT 27.410 10.150 29.235 10.175 ;
        RECT 60.125 6.825 60.565 47.085 ;
        RECT 65.685 43.645 66.125 47.085 ;
        RECT 65.635 43.170 66.175 43.645 ;
        RECT 132.280 38.060 134.385 40.865 ;
        RECT 123.645 26.450 124.025 26.880 ;
        RECT 136.120 26.875 137.120 27.700 ;
        RECT 122.840 26.030 124.025 26.450 ;
        RECT 89.275 25.340 90.255 25.680 ;
        RECT 108.215 20.085 108.595 24.350 ;
        RECT 103.630 19.300 108.595 20.085 ;
        RECT 93.520 13.370 93.970 15.220 ;
        RECT 89.275 13.030 93.970 13.370 ;
        RECT 68.700 10.880 80.265 12.005 ;
        RECT 93.520 10.460 93.970 13.030 ;
        RECT 97.960 13.010 98.415 15.220 ;
        RECT 93.470 9.915 94.020 10.460 ;
        RECT 39.570 5.925 60.565 6.825 ;
        RECT 39.570 3.925 40.470 5.925 ;
        RECT 39.520 3.100 40.520 3.925 ;
        RECT 97.480 3.425 98.485 4.220 ;
        RECT 103.630 4.205 104.415 19.300 ;
        RECT 122.840 14.050 123.260 26.030 ;
        RECT 123.645 25.990 124.025 26.030 ;
        RECT 105.065 10.150 106.690 12.040 ;
        RECT 121.665 7.115 122.425 7.910 ;
        RECT 103.630 3.420 117.780 4.205 ;
        RECT 58.840 3.005 59.840 3.415 ;
        RECT 78.160 1.925 79.160 2.300 ;
      LAYER met4 ;
        RECT 78.810 224.760 78.815 225.290 ;
        RECT 15.030 219.655 15.330 224.760 ;
        RECT 17.790 219.655 18.090 224.760 ;
        RECT 20.550 219.655 20.850 224.760 ;
        RECT 23.310 219.655 23.610 224.760 ;
        RECT 26.070 219.655 26.370 224.760 ;
        RECT 28.830 219.655 29.130 224.760 ;
        RECT 31.590 219.655 31.890 224.760 ;
        RECT 34.350 219.655 34.650 224.760 ;
        RECT 37.110 219.655 37.410 224.760 ;
        RECT 39.870 219.655 40.170 224.760 ;
        RECT 42.630 219.655 42.930 224.760 ;
        RECT 45.390 219.655 45.690 224.760 ;
        RECT 48.150 219.655 48.450 224.760 ;
        RECT 50.910 219.655 51.210 224.760 ;
        RECT 53.670 219.655 53.970 224.760 ;
        RECT 56.430 219.655 56.730 224.760 ;
        RECT 59.190 219.655 59.490 224.760 ;
        RECT 61.950 219.655 62.250 224.760 ;
        RECT 64.710 219.655 65.010 224.760 ;
        RECT 67.470 219.655 67.770 224.760 ;
        RECT 70.230 219.655 70.530 224.760 ;
        RECT 72.990 219.655 73.290 224.760 ;
        RECT 75.750 219.655 76.050 224.760 ;
        RECT 78.510 219.655 78.815 224.760 ;
        RECT 6.000 218.705 78.825 219.655 ;
        RECT 78.510 218.700 78.815 218.705 ;
        RECT 57.615 183.905 87.225 213.515 ;
        RECT 82.510 181.235 85.825 183.905 ;
        RECT 88.580 183.570 89.060 213.850 ;
        RECT 92.095 183.915 121.705 213.525 ;
        RECT 57.610 154.535 87.220 181.235 ;
        RECT 53.005 154.025 87.220 154.535 ;
        RECT 10.225 152.285 12.235 152.290 ;
        RECT 6.000 150.285 12.235 152.285 ;
        RECT 10.225 150.280 12.235 150.285 ;
        RECT 55.340 148.970 56.130 154.025 ;
        RECT 57.610 151.625 87.220 154.025 ;
        RECT 84.040 149.500 87.185 151.625 ;
        RECT 88.575 151.290 89.055 181.570 ;
        RECT 94.125 181.225 97.295 183.915 ;
        RECT 123.060 183.580 123.540 213.860 ;
        RECT 92.090 151.615 121.700 181.225 ;
        RECT 92.140 149.500 95.350 151.615 ;
        RECT 123.055 151.280 123.535 181.560 ;
        RECT 55.335 147.990 56.135 148.970 ;
        RECT 84.040 146.350 95.350 149.500 ;
        RECT 125.435 150.855 127.200 150.860 ;
        RECT 125.435 149.295 142.000 150.855 ;
        RECT 125.435 149.290 127.200 149.295 ;
        RECT 31.175 139.910 35.480 139.920 ;
        RECT 6.000 137.910 35.480 139.910 ;
        RECT 31.175 137.905 35.480 137.910 ;
        RECT 27.495 120.575 27.995 120.580 ;
        RECT 21.825 120.225 28.210 120.575 ;
        RECT 21.825 49.600 22.490 120.225 ;
        RECT 27.495 120.220 27.995 120.225 ;
        RECT 55.540 109.220 56.050 109.730 ;
        RECT 30.840 98.435 31.235 98.440 ;
        RECT 30.040 97.935 31.280 98.435 ;
        RECT 26.360 96.920 26.870 97.315 ;
        RECT 26.365 55.630 26.865 96.920 ;
        RECT 30.040 88.200 30.540 97.935 ;
        RECT 30.840 97.930 31.235 97.935 ;
        RECT 30.040 87.700 32.035 88.200 ;
        RECT 31.705 87.190 32.035 87.700 ;
        RECT 55.545 85.810 56.045 109.220 ;
        RECT 110.340 107.700 110.820 135.480 ;
        RECT 112.175 108.035 139.285 135.145 ;
        RECT 112.175 106.265 115.280 108.035 ;
        RECT 107.010 105.755 115.280 106.265 ;
        RECT 100.630 104.740 101.140 105.250 ;
        RECT 99.070 92.690 99.400 95.200 ;
        RECT 100.635 92.690 101.135 104.740 ;
        RECT 107.010 93.655 107.520 105.755 ;
        RECT 99.070 92.190 101.135 92.690 ;
        RECT 57.150 85.810 57.480 88.320 ;
        RECT 55.545 85.310 57.480 85.810 ;
        RECT 55.545 76.300 56.045 85.310 ;
        RECT 100.635 83.180 101.135 92.190 ;
        RECT 57.150 82.680 101.135 83.180 ;
        RECT 57.150 80.170 57.480 82.680 ;
        RECT 110.340 76.770 110.820 104.550 ;
        RECT 112.175 104.215 115.280 105.755 ;
        RECT 112.175 77.105 139.285 104.215 ;
        RECT 55.545 75.800 99.400 76.300 ;
        RECT 99.070 73.910 99.400 75.800 ;
        RECT 47.955 72.320 110.635 72.370 ;
        RECT 47.955 69.905 142.000 72.320 ;
        RECT 47.955 65.300 50.625 69.905 ;
        RECT 60.385 69.870 64.470 69.905 ;
        RECT 107.625 69.895 110.275 69.905 ;
        RECT 107.625 69.890 110.270 69.895 ;
        RECT 47.950 64.630 50.630 65.300 ;
        RECT 61.745 60.510 64.470 69.870 ;
        RECT 61.740 59.625 64.475 60.510 ;
        RECT 26.360 55.260 26.870 55.630 ;
        RECT 30.845 52.415 40.420 52.815 ;
        RECT 30.845 51.630 31.175 52.415 ;
        RECT 21.820 49.085 22.495 49.600 ;
        RECT 19.620 48.335 20.295 48.845 ;
        RECT 14.335 42.645 16.335 42.650 ;
        RECT 6.000 40.645 16.335 42.645 ;
        RECT 14.335 40.640 16.335 40.645 ;
        RECT 14.950 12.010 16.785 12.015 ;
        RECT 6.000 10.175 16.785 12.010 ;
        RECT 14.950 10.170 16.785 10.175 ;
        RECT 19.625 7.805 20.290 48.335 ;
        RECT 39.920 47.605 40.420 52.415 ;
        RECT 45.175 50.835 45.505 51.525 ;
        RECT 45.175 50.515 54.275 50.835 ;
        RECT 38.215 47.105 40.420 47.605 ;
        RECT 38.215 43.700 38.545 47.105 ;
        RECT 52.525 45.410 52.855 46.100 ;
        RECT 53.955 45.410 54.275 50.515 ;
        RECT 52.525 45.090 54.275 45.410 ;
        RECT 38.210 43.370 38.550 43.700 ;
        RECT 52.525 43.645 52.855 45.090 ;
        RECT 65.680 43.645 66.130 43.650 ;
        RECT 52.525 43.170 66.130 43.645 ;
        RECT 30.800 41.940 31.225 41.945 ;
        RECT 27.245 41.610 43.375 41.940 ;
        RECT 30.800 41.605 31.225 41.610 ;
        RECT 43.045 37.745 43.375 41.610 ;
        RECT 52.525 41.435 52.855 43.170 ;
        RECT 65.680 43.165 66.130 43.170 ;
        RECT 25.485 37.415 43.375 37.745 ;
        RECT 25.485 34.780 25.815 37.415 ;
        RECT 25.485 34.450 27.575 34.780 ;
        RECT 43.045 34.320 43.375 37.415 ;
        RECT 45.560 40.530 46.370 40.860 ;
        RECT 132.325 40.840 134.340 40.845 ;
        RECT 45.560 34.320 45.880 40.530 ;
        RECT 132.325 38.085 142.000 40.840 ;
        RECT 132.325 38.080 134.340 38.085 ;
        RECT 43.045 34.000 45.880 34.320 ;
        RECT 43.045 31.200 43.375 34.000 ;
        RECT 41.810 30.870 43.375 31.200 ;
        RECT 136.165 26.895 137.075 27.680 ;
        RECT 89.320 25.345 98.375 25.675 ;
        RECT 97.995 13.045 98.375 25.345 ;
        RECT 98.005 13.030 98.370 13.045 ;
        RECT 105.110 12.010 106.645 12.020 ;
        RECT 27.405 10.175 106.675 12.010 ;
        RECT 105.110 10.170 106.645 10.175 ;
        RECT 121.710 7.805 122.380 7.890 ;
        RECT 19.625 7.140 122.380 7.805 ;
        RECT 121.710 7.135 122.380 7.140 ;
        RECT 121.715 7.090 122.380 7.135 ;
        RECT 97.530 4.200 98.435 4.515 ;
        RECT 39.565 3.095 40.475 3.930 ;
        RECT 97.525 3.445 98.440 4.200 ;
        RECT 39.570 1.000 40.470 3.095 ;
        RECT 58.885 3.000 59.795 3.395 ;
        RECT 58.890 1.000 59.790 3.000 ;
        RECT 78.205 1.920 79.115 2.280 ;
        RECT 78.210 1.000 79.110 1.920 ;
        RECT 97.530 1.000 98.435 3.445 ;
        RECT 116.845 3.415 117.755 4.210 ;
        RECT 116.850 1.000 117.750 3.415 ;
        RECT 136.170 1.000 137.070 26.895 ;
        RECT 98.430 0.940 98.435 1.000 ;
  END
END tt_um_DalinEM_asic
END LIBRARY

